netcdf CFS-atmos-northPacific-rain-2017 {
dimensions:
	lat = 344 ;
	lon = 588 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double rain(rain_time, lat, lon) ;
		rain:missing_value = -1.e+34 ;
		rain:_FillValue = -1.e+34 ;
		rain:time = "rain_time" ;
		rain:coordinates = "lon lat" ;
		rain:long_name = "rainfall" ;
		rain:history = "From roms-cfs-atmos-rain-2017" ;
	double rain_time(rain_time) ;
		rain_time:units = "day since 1900-01-01 00:00:00" ;
		rain_time:time_origin = "01-JAN-1900 00:00:00" ;
		rain_time:axis = "T" ;
		rain_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:20:44 2022: ncks -F -O -d rain_time,3,1462 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2017/roms-cfs-atmos-rain-2017.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-rain-2017.nc\n",
			"Mon Sep 17 12:11:07 2018: Time overhang added\n",
			"Mon Sep 17 12:10:59 2018: ncrcat /tmp/tp48d98b7d_b445_4ffb_8f68_15e50fd01480.nc frc/roms-cfs-atmos-rain-2017.nc /tmp/tp277bcd3b_1a47_444f_96fd_e2302d4973a9.nc /tmp/tpab1718f1_3314_44d2_9bd0_895fc4b0957d.nc\n",
			"Mon Sep 17 12:10:59 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2017.nc /tmp/tp48d98b7d_b445_4ffb_8f68_15e50fd01480.nc\n",
			"FERRET V7.4  10-Aug-18" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
