netcdf CFS-atmos-northPacific-rain-1997 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:40 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1997/roms-cfs-atmos-rain-1997.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1997/CFS-atmos-northPacific-rain-1997.nc\n",
			"Mon Sep 10 13:49:55 2018: Time overhang added\n",
			"Mon Sep 10 13:49:51 2018: ncrcat /tmp/tpf2ebb8e9_57fa_4b34_bf13_3ab34201e6c7.nc frc/roms-cfs-atmos-rain-1997.nc /tmp/tp01bfe9ae_b6ee_41fa_b826_821f04ac2073.nc /tmp/tpa6f369af_2acc_47af_8779_ab8a67af037f.nc\n",
			"Mon Sep 10 13:49:51 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-1997.nc /tmp/tpf2ebb8e9_57fa_4b34_bf13_3ab34201e6c7.nc\n",
			"Thu Sep  6 10:10:32 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1997_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-1997.nc\n",
			"04-Oct-2017 17:43:50: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
