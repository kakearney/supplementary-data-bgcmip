netcdf INIbgc_BIO_COBALT_NEP {
dimensions:
	xi_rho = 226 ;
	eta_rho = 642 ;
	s_rho = 30 ;
	ocean_time = UNLIMITED ; // (1 currently)
variables:
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 1900-01-01 00:00:00" ;
		ocean_time:calendar = "standard" ;
	double nsm(ocean_time, s_rho, eta_rho, xi_rho) ;
		nsm:long_name = "Small Phytoplankton Nitrogen" ;
		nsm:unit = "mol/kg" ;
		nsm:time = "ocean_time" ;
		nsm:_FillValue = 1.e+36 ;
	double nlg(ocean_time, s_rho, eta_rho, xi_rho) ;
		nlg:long_name = "Large Phytoplankton Nitrogen" ;
		nlg:unit = "mol/kg" ;
		nlg:time = "ocean_time" ;
		nlg:_FillValue = 1.e+36 ;
	double ndi(ocean_time, s_rho, eta_rho, xi_rho) ;
		ndi:long_name = "Diazotroph Nitrogen" ;
		ndi:unit = "mol/kg" ;
		ndi:time = "ocean_time" ;
		ndi:_FillValue = 1.e+36 ;
	double nsmz(ocean_time, s_rho, eta_rho, xi_rho) ;
		nsmz:long_name = "Small Zooplankton Nitrogen" ;
		nsmz:unit = "mol/kg" ;
		nsmz:time = "ocean_time" ;
		nsmz:_FillValue = 1.e+36 ;
	double nmdz(ocean_time, s_rho, eta_rho, xi_rho) ;
		nmdz:long_name = "Medium-sized zooplankton Nitrogen" ;
		nmdz:unit = "mol/kg" ;
		nmdz:time = "ocean_time" ;
		nmdz:_FillValue = 1.e+36 ;
	double nlgz(ocean_time, s_rho, eta_rho, xi_rho) ;
		nlgz:long_name = "large Zooplankton Nitrogen" ;
		nlgz:unit = "mol/kg" ;
		nlgz:time = "ocean_time" ;
		nlgz:_FillValue = 1.e+36 ;
	double ldon(ocean_time, s_rho, eta_rho, xi_rho) ;
		ldon:long_name = "labile DON" ;
		ldon:unit = "mol/kg" ;
		ldon:time = "ocean_time" ;
		ldon:_FillValue = 1.e+36 ;
	double sldon(ocean_time, s_rho, eta_rho, xi_rho) ;
		sldon:long_name = "Semilabile DON" ;
		sldon:unit = "mol/kg" ;
		sldon:time = "ocean_time" ;
		sldon:_FillValue = 1.e+36 ;
	double srdon(ocean_time, s_rho, eta_rho, xi_rho) ;
		srdon:long_name = "Semi-Refractory DON" ;
		srdon:unit = "mol/kg" ;
		srdon:time = "ocean_time" ;
		srdon:_FillValue = 1.e+36 ;
	double nbact(ocean_time, s_rho, eta_rho, xi_rho) ;
		nbact:long_name = "bacterial" ;
		nbact:unit = "mol/kg" ;
		nbact:time = "ocean_time" ;
		nbact:_FillValue = 1.e+36 ;
	double nh4(ocean_time, s_rho, eta_rho, xi_rho) ;
		nh4:long_name = "Ammonia" ;
		nh4:unit = "mol/kg" ;
		nh4:time = "ocean_time" ;
		nh4:_FillValue = 1.e+36 ;
	double no3(ocean_time, s_rho, eta_rho, xi_rho) ;
		no3:long_name = "Nitrate" ;
		no3:unit = "mol/kg" ;
		no3:time = "ocean_time" ;
		no3:_FillValue = 1.e+36 ;
	double ndet(ocean_time, s_rho, eta_rho, xi_rho) ;
		ndet:long_name = "ndet" ;
		ndet:unit = "mol/kg" ;
		ndet:time = "ocean_time" ;
		ndet:_FillValue = 1.e+36 ;
	double sio4(ocean_time, s_rho, eta_rho, xi_rho) ;
		sio4:long_name = "Silicate" ;
		sio4:unit = "mol/kg" ;
		sio4:time = "ocean_time" ;
		sio4:_FillValue = 1.e+36 ;
	double silg(ocean_time, s_rho, eta_rho, xi_rho) ;
		silg:long_name = "Large Phytoplankton Silicon" ;
		silg:unit = "mol/kg" ;
		silg:time = "ocean_time" ;
		silg:_FillValue = 1.e+36 ;
	double sidet(ocean_time, s_rho, eta_rho, xi_rho) ;
		sidet:long_name = "Detrital Silicon" ;
		sidet:unit = "mol/kg" ;
		sidet:time = "ocean_time" ;
		sidet:_FillValue = 1.e+36 ;
	double cadet_calc(ocean_time, s_rho, eta_rho, xi_rho) ;
		cadet_calc:long_name = "Detrital CaCO3" ;
		cadet_calc:unit = "mol/kg" ;
		cadet_calc:time = "ocean_time" ;
		cadet_calc:_FillValue = 1.e+36 ;
	double cadet_arag(ocean_time, s_rho, eta_rho, xi_rho) ;
		cadet_arag:long_name = "Detrital CaCO3" ;
		cadet_arag:unit = "mol/kg" ;
		cadet_arag:time = "ocean_time" ;
		cadet_arag:_FillValue = 1.e+36 ;
	double lith(ocean_time, s_rho, eta_rho, xi_rho) ;
		lith:long_name = "Lithogenic Aluminosilicate" ;
		lith:unit = "g/kg" ;
		lith:time = "ocean_time" ;
		lith:_FillValue = 1.e+36 ;
	double lithdet(ocean_time, s_rho, eta_rho, xi_rho) ;
		lithdet:long_name = "lithdet" ;
		lithdet:unit = "g/kg" ;
		lithdet:time = "ocean_time" ;
		lithdet:_FillValue = 1.e+36 ;
	double po4(ocean_time, s_rho, eta_rho, xi_rho) ;
		po4:long_name = "Phosphate" ;
		po4:unit = "mol/kg" ;
		po4:time = "ocean_time" ;
		po4:_FillValue = 1.e+36 ;
	double ldop(ocean_time, s_rho, eta_rho, xi_rho) ;
		ldop:long_name = "labile DOP" ;
		ldop:unit = "mol/kg" ;
		ldop:time = "ocean_time" ;
		ldop:_FillValue = 1.e+36 ;
	double sldop(ocean_time, s_rho, eta_rho, xi_rho) ;
		sldop:long_name = "Semilabile DOP" ;
		sldop:unit = "mol/kg" ;
		sldop:time = "ocean_time" ;
		sldop:_FillValue = 1.e+36 ;
	double srdop(ocean_time, s_rho, eta_rho, xi_rho) ;
		srdop:long_name = "Semi-Refractory DOP" ;
		srdop:unit = "mol/kg" ;
		srdop:time = "ocean_time" ;
		srdop:_FillValue = 1.e+36 ;
	double pdet(ocean_time, s_rho, eta_rho, xi_rho) ;
		pdet:long_name = "Detrital Phosphorus" ;
		pdet:unit = "mol/kg" ;
		pdet:time = "ocean_time" ;
		pdet:_FillValue = 1.e+36 ;
	double fesm(ocean_time, s_rho, eta_rho, xi_rho) ;
		fesm:long_name = "Small Phytoplankton Iron" ;
		fesm:unit = "mol/kg" ;
		fesm:time = "ocean_time" ;
		fesm:_FillValue = 1.e+36 ;
	double fedi(ocean_time, s_rho, eta_rho, xi_rho) ;
		fedi:long_name = "Diazotroph Iron" ;
		fedi:unit = "mol/kg" ;
		fedi:time = "ocean_time" ;
		fedi:_FillValue = 1.e+36 ;
	double felg(ocean_time, s_rho, eta_rho, xi_rho) ;
		felg:long_name = "Large Phytoplankton Iron" ;
		felg:unit = "mol/kg" ;
		felg:time = "ocean_time" ;
		felg:_FillValue = 1.e+36 ;
	double fed(ocean_time, s_rho, eta_rho, xi_rho) ;
		fed:long_name = "Dissolved Iron" ;
		fed:unit = "mol/kg" ;
		fed:time = "ocean_time" ;
		fed:_FillValue = 1.e+36 ;
	double fedet(ocean_time, s_rho, eta_rho, xi_rho) ;
		fedet:long_name = "Detrital Iron" ;
		fedet:unit = "mol/kg" ;
		fedet:time = "ocean_time" ;
		fedet:_FillValue = 1.e+36 ;
	double o2(ocean_time, s_rho, eta_rho, xi_rho) ;
		o2:long_name = "Oxygen" ;
		o2:unit = "mol/kg" ;
		o2:time = "ocean_time" ;
		o2:_FillValue = 1.e+36 ;
	double dic(ocean_time, s_rho, eta_rho, xi_rho) ;
		dic:long_name = "Dissolved Inorganic Carbon" ;
		dic:unit = "mol/kg" ;
		dic:time = "ocean_time" ;
		dic:_FillValue = 1.e+36 ;
	double alk(ocean_time, s_rho, eta_rho, xi_rho) ;
		alk:long_name = "Alkalinity" ;
		alk:unit = "mol/kg" ;
		alk:time = "ocean_time" ;
		alk:_FillValue = 1.e+36 ;
	double nmd(ocean_time, s_rho, eta_rho, xi_rho) ;
		nmd:long_name = "Medium Phytoplankton Nitrogen" ;
		nmd:unit = "mol/kg" ;
		nmd:time = "ocean_time" ;
		nmd:_FillValue = 1.e+36 ;
	double simd(ocean_time, s_rho, eta_rho, xi_rho) ;
		simd:long_name = "Medium Phytoplankton Silicon" ;
		simd:unit = "mol/kg" ;
		simd:time = "ocean_time" ;
		simd:_FillValue = 1.e+36 ;
	double femd(ocean_time, s_rho, eta_rho, xi_rho) ;
		femd:long_name = "Medium Phytoplankton Iron" ;
		femd:unit = "mol/kg" ;
		femd:time = "ocean_time" ;
		femd:_FillValue = 1.e+36 ;
	double cased(ocean_time, s_rho, eta_rho, xi_rho) ;
		cased:long_name = "Sediment CaCO3" ;
		cased:unit = "mol m-3" ;
		cased:time = "ocean_time" ;
		cased:_FillValue = 1.e+36 ;
	double cadet_arag_btf(ocean_time, eta_rho, xi_rho) ;
		cadet_arag_btf:long_name = "aragonite flux to Sediments" ;
		cadet_arag_btf:unit = "mol m-2 s-1" ;
		cadet_arag_btf:time = "ocean_time" ;
		cadet_arag_btf:_FillValue = 1.e+36 ;
	double cadet_calc_btf(ocean_time, eta_rho, xi_rho) ;
		cadet_calc_btf:long_name = "calcite flux to Sediments" ;
		cadet_calc_btf:unit = "mol m-2 s-1" ;
		cadet_calc_btf:time = "ocean_time" ;
		cadet_calc_btf:_FillValue = 1.e+36 ;
	double ndet_btf(ocean_time, eta_rho, xi_rho) ;
		ndet_btf:long_name = "N flux to Sediments" ;
		ndet_btf:unit = "mol m-2 s-1" ;
		ndet_btf:time = "ocean_time" ;
		ndet_btf:_FillValue = 1.e+36 ;
	double pdet_btf(ocean_time, eta_rho, xi_rho) ;
		pdet_btf:long_name = "P flux to Sediments" ;
		pdet_btf:unit = "mol m-2 s-1" ;
		pdet_btf:time = "ocean_time" ;
		pdet_btf:_FillValue = 1.e+36 ;
	double sidet_btf(ocean_time, eta_rho, xi_rho) ;
		sidet_btf:long_name = "SiO2 flux to Sediments" ;
		sidet_btf:unit = "mol m-2 s-1" ;
		sidet_btf:time = "ocean_time" ;
		sidet_btf:_FillValue = 1.e+36 ;
	double chl(ocean_time, s_rho, eta_rho, xi_rho) ;
		chl:long_name = "Chlorophyll" ;
		chl:unit = "ug/kg" ;
		chl:time = "ocean_time" ;
		chl:_FillValue = 1.e+36 ;
	double irr_mem(ocean_time, s_rho, eta_rho, xi_rho) ;
		irr_mem:long_name = "Irradiance memory" ;
		irr_mem:unit = "Watts/m^2" ;
		irr_mem:time = "ocean_time" ;
		irr_mem:_FillValue = 1.e+36 ;
	double htotal(ocean_time, s_rho, eta_rho, xi_rho) ;
		htotal:long_name = "H+ ion concentration" ;
		htotal:unit = "mol/kg" ;
		htotal:time = "ocean_time" ;
		htotal:_FillValue = 1.e+36 ;
	double co3_ion(ocean_time, s_rho, eta_rho, xi_rho) ;
		co3_ion:long_name = "Carbonate ion" ;
		co3_ion:unit = "mol/kg" ;
		co3_ion:time = "ocean_time" ;
		co3_ion:_FillValue = 1.e+36 ;
	double mu_mem_sm(ocean_time, s_rho, eta_rho, xi_rho) ;
		mu_mem_sm:long_name = "Aggreg memory small phyto" ;
		mu_mem_sm:time = "ocean_time" ;
		mu_mem_sm:_FillValue = 1.e+36 ;
	double mu_mem_di(ocean_time, s_rho, eta_rho, xi_rho) ;
		mu_mem_di:long_name = "Aggreg memory diatoms" ;
		mu_mem_di:time = "ocean_time" ;
		mu_mem_di:_FillValue = 1.e+36 ;
	double mu_mem_lg(ocean_time, s_rho, eta_rho, xi_rho) ;
		mu_mem_lg:long_name = "Aggreg memory large phyto" ;
		mu_mem_lg:time = "ocean_time" ;
		mu_mem_lg:_FillValue = 1.e+36 ;
	double mu_mem_md(ocean_time, s_rho, eta_rho, xi_rho) ;
		mu_mem_md:long_name = "Aggreg memory medium phyto" ;
		mu_mem_md:time = "ocean_time" ;
		mu_mem_md:_FillValue = 1.e+36 ;

// global attributes:
		:type = "INITIALIZATION file" ;
		:history = "Wed Jan 25 11:27:16 2023: BGC data added: NO3, PO4, Alk, TIC, O2, SiO4: GLODAPv2.2016b Mapped Climatologies; Fe: Huang et al., 2022 climatology + GOANPZ analytical; Hfree, CO3: GLODAPv2 + CO2sys; producers/consumers: seed value; others: 0\n",
			"Wed Jan 25 11:27:11 2023: File schema created via ini_schema.m" ;
}
