netcdf CFS-atmos-northPacific-rain-2015 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:53:05 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2015/roms-cfs-atmos-rain-2015.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-rain-2015.nc\n",
			"Mon Sep 10 14:03:02 2018: Time overhang added\n",
			"Mon Sep 10 14:02:55 2018: ncrcat /tmp/tp9db026a0_fad3_441e_8884_42b349012569.nc frc/roms-cfs-atmos-rain-2015.nc /tmp/tp3740aef5_19ce_4e34_b4c1_3dbaa1974e30.nc /tmp/tpe5af171d_0280_47cd_84ee_ee3f464369d7.nc\n",
			"Mon Sep 10 14:02:54 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2015.nc /tmp/tp9db026a0_fad3_441e_8884_42b349012569.nc\n",
			"Thu Sep  6 13:51:10 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2015_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2015.nc\n",
			"04-Oct-2017 18:32:06: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
