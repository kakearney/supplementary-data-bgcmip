netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2021 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 17:02:43 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:59:51 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2021/CFS-ocean-NEP-N30-bryocn-2021.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2021/CFS-ocean-ESPER-NEP-N30-brycarbon-2021.nc\n",
			"Fri Jan 13 10:35:10 2023: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad73.nc <>/final/2021/CFS-ocean-NEP-N30-bryocn-2021.nc\n",
			"Fri Jan 13 10:32:47 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad01.nc\n",
			"Fri Jan 13 10:32:47 2023: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad01.nc\n",
			"Fri Jan 13 10:32:46 2023: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2021010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2021pentad01.nc\n",
			"Thu Jan 12 22:12:12 2023: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
