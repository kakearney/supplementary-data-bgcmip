netcdf CFS-atmos-northPacific-Qair-2004 {
dimensions:
	qair_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:50:41 2022: ncks -F -O -d qair_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2004/roms-cfs-atmos-Qair-2004.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2004/CFS-atmos-northPacific-Qair-2004.nc\n",
			"Mon Sep 10 13:35:22 2018: Time overhang added\n",
			"Mon Sep 10 13:35:18 2018: ncrcat /tmp/tpd29fbe7c_1818_4cd3_a3c8_00c1bb0b7278.nc frc/roms-cfs-atmos-Qair-2004.nc /tmp/tpb96c5eb6_4626_4e64_aebf_180ebf8767e2.nc /tmp/tp190d73ef_c129_41b1_956d_7664171ba72b.nc\n",
			"Mon Sep 10 13:35:18 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2004.nc /tmp/tpd29fbe7c_1818_4cd3_a3c8_00c1bb0b7278.nc\n",
			"Thu Sep  6 11:11:33 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2004.nc\n",
			"Thu Sep  6 11:10:45 2018: ncks -O -F -d air_time,2,1465 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2004_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2004.nc\n",
			"04-Oct-2017 17:59:35: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
