netcdf CFS-atmos-northPacific-rain-2002 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:41 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2002/roms-cfs-atmos-rain-2002.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2002/CFS-atmos-northPacific-rain-2002.nc\n",
			"Mon Sep 10 13:50:24 2018: Time overhang added\n",
			"Mon Sep 10 13:50:20 2018: ncrcat /tmp/tp8b5e7e8e_ad7d_4b7b_b9f9_211f69d3e0c4.nc frc/roms-cfs-atmos-rain-2002.nc /tmp/tp8b01e57f_5e32_43f2_be2c_6759f4faccff.nc /tmp/tp7c1359d0_07e5_4628_9cc4_5122fd16a75c.nc\n",
			"Mon Sep 10 13:50:20 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2002.nc /tmp/tp8b5e7e8e_ad7d_4b7b_b9f9_211f69d3e0c4.nc\n",
			"Thu Sep  6 10:55:36 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2002_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2002.nc\n",
			"04-Oct-2017 17:56:46: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
