netcdf CFS-atmos-northPacific-Qair-1985 {
dimensions:
	qair_time = UNLIMITED ; // (1459 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:missing_value = -1.e+34 ;
		Qair:_FillValue = -1.e+34 ;
		Qair:time = "qair_time" ;
		Qair:coordinates = "lon lat" ;
		Qair:height_above_ground = 2.f ;
		Qair:long_name = "specific humidity" ;
		Qair:history = "From roms-cfs-atmos-Qair-1985" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double qair_time(qair_time) ;
		qair_time:units = "day since 1900-01-01 00:00:00" ;
		qair_time:time_origin = "01-JAN-1900 00:00:00" ;
		qair_time:axis = "T" ;
		qair_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:18:44 2022: ncks -F -O -d qair_time,2,1460 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1985/roms-cfs-atmos-Qair-1985.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1985/CFS-atmos-northPacific-Qair-1985.nc\n",
			"Wed Nov 20 13:46:15 2019: Time overhang added to end\n",
			"Wed Nov 20 13:46:10 2019: ncrcat /gscratch/bumblereem/bering10k/input/hindcast_cfs/1985/roms-cfs-atmos-Qair-1985.nc /tmp/tpb47b3940_2c7c_46e3_b70e_79404be43347.nc /tmp/tp0f3ec65b_2b83_4e6b_87d0_65a871b8a279.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
