netcdf CFS-atmos-northPacific-Uwind-1998 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:45:41 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1998/roms-cfs-atmos-Uwind-1998.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1998/CFS-atmos-northPacific-Uwind-1998.nc\n",
			"Mon Sep 10 13:40:40 2018: Time overhang added\n",
			"Mon Sep 10 13:40:37 2018: ncrcat /tmp/tp98ee256f_f22a_4934_9769_2020a6477e44.nc frc/roms-cfs-atmos-Uwind-1998.nc /tmp/tp9317cb7b_eb8b_422b_96de_8e6b5880c78f.nc /tmp/tp0d60e0c4_ce46_4afd_b4b7_101a037e3dae.nc\n",
			"Mon Sep 10 13:40:37 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-1998.nc /tmp/tp98ee256f_f22a_4934_9769_2020a6477e44.nc\n",
			"Thu Sep  6 10:18:31 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1998_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-1998.nc\n",
			"04-Oct-2017 17:45:35: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
