netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-1994 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 14:45:48 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 14:42:53 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1994/CFS-ocean-NEP-N30-bryocn-1994.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1994/CFS-ocean-ESPER-NEP-N30-brycarbon-1994.nc\n",
			"Thu Dec 15 10:03:37 2022: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad73.nc <>/final/1994/CFS-ocean-NEP-N30-bryocn-1994.nc\n",
			"Thu Dec 15 10:02:52 2022: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad01.nc\n",
			"Thu Dec 15 10:02:52 2022: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1994010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1994pentad01.nc\n",
			"Wed Dec 14 19:34:47 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
