netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-1995 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 14:48:02 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 14:46:16 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1995/CFS-ocean-Bering10K-N30-bryocn-1995.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1995/CFS-ocean-ESPER-Bering10K-N30-brycarbon-1995.nc\n",
			"Fri Dec 16 01:03:48 2022: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad73.nc <>/final/1995/CFS-ocean-Bering10K-N30-bryocn-1995.nc\n",
			"Fri Dec 16 01:03:07 2022: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad01.nc\n",
			"Fri Dec 16 01:03:06 2022: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1995010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1995pentad01.nc\n",
			"Thu Dec 15 10:04:50 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
