netcdf CFS-atmos-northPacific-swrad-1997 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:45 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1997/roms-cfs-atmos-swrad-1997.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1997/CFS-atmos-northPacific-swrad-1997.nc\n",
			"Mon Sep 10 14:03:44 2018: Time overhang added\n",
			"Mon Sep 10 14:03:43 2018: ncrcat /tmp/tpe692353f_70c6_4ab6_ac80_a631d690d8ad.nc frc/roms-cfs-atmos-swrad-1997.nc /tmp/tpdd76de10_64d6_4f1d_842c_c2953edd10d5.nc /tmp/tp0520f2e6_53ce_4783_8acf_3e4f162f286e.nc\n",
			"Mon Sep 10 14:03:43 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-1997.nc /tmp/tpe692353f_70c6_4ab6_ac80_a631d690d8ad.nc\n",
			"Thu Sep  6 10:11:06 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1997_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-1997.nc\n",
			"04-Oct-2017 17:43:00: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
