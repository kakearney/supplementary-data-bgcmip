netcdf CFS-atmos-northPacific-Tair-2020 {
dimensions:
	tair_time = UNLIMITED ; // (1448 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:missing_value = -1.e+34 ;
		Tair:_FillValue = -1.e+34 ;
		Tair:time = "tair_time" ;
		Tair:coordinates = "lon lat" ;
		Tair:height_above_ground = 2.f ;
		Tair:long_name = "surface air temperature" ;
		Tair:history = "From roms-cfs-atmos-Tair-2020" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double tair_time(tair_time) ;
		tair_time:units = "day since 1900-01-01 00:00:00" ;
		tair_time:time_origin = "01-JAN-1900 00:00:00" ;
		tair_time:axis = "T" ;
		tair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:52:57 2022: ncks -F -O -d tair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Tair-2020.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Tair-2020.nc\n",
			"Wed Jan 27 10:11:17 2021: Time overhang added to both ends\n",
			"Wed Jan 27 10:11:08 2021: ncrcat /tmp/tpa0614985_6185_4a21_94e2_b6298e48a457.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Tair-2020.nc /tmp/tp02fbe600_7679_4239_9e78_e7c1562a4072.nc /tmp/tp723a8f7c_b633_40d8_b1e5_17db87fbfa99.nc\n",
			"Wed Jan 27 10:11:07 2021: ncks -F -d tair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Tair-2020.nc /tmp/tpa0614985_6185_4a21_94e2_b6298e48a457.nc\n",
			"FERRET V7.6  26-Jan-21" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
