netcdf CFS-atmos-northPacific-Tair-2013 {
dimensions:
	tair_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:22:04 2022: ncks -F -O -d tair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2013/roms-cfs-atmos-Tair-2013.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Tair-2013.nc\n",
			"Mon Sep 10 13:39:23 2018: Time overhang added\n",
			"Mon Sep 10 13:39:15 2018: ncrcat /tmp/tp3c7247c6_5ab4_41bf_9aad_6e92433d153a.nc frc/roms-cfs-atmos-Tair-2013.nc /tmp/tp98bdf21d_c6a4_45a5_800f_7883ce9455b8.nc /tmp/tp3f01f974_4920_4ac8_adc4_3a712e5d8847.nc\n",
			"Mon Sep 10 13:39:14 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2013.nc /tmp/tp3c7247c6_5ab4_41bf_9aad_6e92433d153a.nc\n",
			"Thu Sep  6 12:56:13 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2013.nc\n",
			"Thu Sep  6 12:54:19 2018: ncks -O -F -d air_time,2,1449 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2013_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2013.nc\n",
			"04-Oct-2017 18:21:22: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
