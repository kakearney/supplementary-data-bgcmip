netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-1990 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 14:22:50 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 14:21:06 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1990/CFS-ocean-ESPER-Bering10K-N30-brycarbon-1990.nc\n",
			"Mon Dec 12 10:29:38 2022: ncrcat -O <>/final/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad73.nc <>/final/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc\n",
			"Fri Dec  9 16:24:34 2022: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad01.nc <>/final/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc\n",
			"Fri Dec  9 16:24:34 2022: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad01.nc\n",
			"Fri Dec  9 16:24:34 2022: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad01.nc\n",
			"Fri Dec 09 16:09:28 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
