netcdf CFS-atmos-northPacific-Pair-1989 {
dimensions:
	pair_time = UNLIMITED ; // (1459 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:missing_value = -1.e+34 ;
		Pair:_FillValue = -1.e+34 ;
		Pair:time = "pair_time" ;
		Pair:coordinates = "lon lat" ;
		Pair:long_name = "atmos pressure" ;
		Pair:history = "From roms-cfs-atmos-Pair-1989" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double pair_time(pair_time) ;
		pair_time:units = "day since 1900-01-01 00:00:00" ;
		pair_time:time_origin = "01-JAN-1900 00:00:00" ;
		pair_time:axis = "T" ;
		pair_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:22:23 2022: ncks -F -O -d pair_time,2,1460 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1989/roms-cfs-atmos-Pair-1989.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1989/CFS-atmos-northPacific-Pair-1989.nc\n",
			"Wed Nov 20 13:54:26 2019: Time overhang added to end\n",
			"Wed Nov 20 13:54:21 2019: ncrcat /gscratch/bumblereem/bering10k/input/hindcast_cfs/1989/roms-cfs-atmos-Pair-1989.nc /tmp/tp59eb7751_3c5c_4066_927b_aaa7e16a1570.nc /tmp/tp7b8c80c3_1426_4ee5_9bcb_6aead7835484.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
