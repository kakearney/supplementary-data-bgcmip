netcdf CFS-atmos-northPacific-Qair-1997 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:08 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1997/roms-cfs-atmos-Qair-1997.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1997/CFS-atmos-northPacific-Qair-1997.nc\n",
			"Mon Sep 10 13:34:43 2018: Time overhang added\n",
			"Mon Sep 10 13:34:40 2018: ncrcat /tmp/tp15aa0c25_ebae_4db8_a246_ba30fc056dfb.nc frc/roms-cfs-atmos-Qair-1997.nc /tmp/tp52b631aa_e566_48d1_b98a_e9eb6f32f56f.nc /tmp/tp9a149597_ee0b_45ab_b46d_df6a37571cf1.nc\n",
			"Mon Sep 10 13:34:39 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-1997.nc /tmp/tp15aa0c25_ebae_4db8_a246_ba30fc056dfb.nc\n",
			"Thu Sep  6 10:09:05 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-1997.nc\n",
			"Thu Sep  6 10:08:19 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1997_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-1997.nc\n",
			"04-Oct-2017 17:41:45: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
