netcdf CFS-atmos-northPacific-Qair-2003 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:56 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2003/roms-cfs-atmos-Qair-2003.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2003/CFS-atmos-northPacific-Qair-2003.nc\n",
			"Mon Sep 10 13:35:16 2018: Time overhang added\n",
			"Mon Sep 10 13:35:13 2018: ncrcat /tmp/tpcff5ccbf_0281_4f14_94c5_cf8b2e789798.nc frc/roms-cfs-atmos-Qair-2003.nc /tmp/tpe7bb3a45_3ba2_4916_8557_0ad0856a9353.nc /tmp/tp581c9e32_1d62_47fc_9974_57b14012fc26.nc\n",
			"Mon Sep 10 13:35:13 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2003.nc /tmp/tpcff5ccbf_0281_4f14_94c5_cf8b2e789798.nc\n",
			"Thu Sep  6 11:03:15 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2003.nc\n",
			"Thu Sep  6 11:02:18 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2003_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2003.nc\n",
			"04-Oct-2017 17:57:09: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
