netcdf CFS-atmos-northPacific-Qair-2011 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:03:04 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2011/roms-cfs-atmos-Qair-2011.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Qair-2011.nc\n",
			"Thu Sep 13 10:47:46 2018: Time overhang added\n",
			"Thu Sep 13 10:47:39 2018: ncrcat /tmp/tp78095084_35b5_4107_967b_39a2676991ab.nc frc/roms-cfs-atmos-Qair-2011.nc /tmp/tp61962063_1407_48a5_bb57_0661571eb0d0.nc /tmp/tp1ea8e7cc_58ef_413e_be46_837cbcaf3a5c.nc\n",
			"Thu Sep 13 10:47:38 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2011.nc /tmp/tp78095084_35b5_4107_967b_39a2676991ab.nc\n",
			"Thu Sep 13 10:42:39 2018: ncrename -d air_time,qair_time -v air_time,qair_time ./frc/roms-cfs-atmos-Qair-2011.nc\n",
			"Thu Sep 13 10:42:29 2018: ncks -O -F -d air_time,2,1461 -v Qair ./frc/Old/corecfs_2011_air.nc ./frc/roms-cfs-atmos-Qair-2011.nc\n",
			"04-Oct-2017 18:13:26: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
