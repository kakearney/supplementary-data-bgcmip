netcdf CFS-atmos-northPacific-Tair-1998 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:45:34 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1998/roms-cfs-atmos-Tair-1998.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1998/CFS-atmos-northPacific-Tair-1998.nc\n",
			"Mon Sep 10 13:37:44 2018: Time overhang added\n",
			"Mon Sep 10 13:37:40 2018: ncrcat /tmp/tpf18180b2_3d0d_486b_a636_83e837a58798.nc frc/roms-cfs-atmos-Tair-1998.nc /tmp/tp063c13d4_32d9_443a_8c3c_588ce5c603d6.nc /tmp/tpfa38f7d1_f640_462a_9708_f2e48c66540f.nc\n",
			"Mon Sep 10 13:37:40 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-1998.nc /tmp/tpf18180b2_3d0d_486b_a636_83e837a58798.nc\n",
			"Thu Sep  6 10:15:16 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1998.nc\n",
			"Thu Sep  6 10:14:18 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1998_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1998.nc\n",
			"04-Oct-2017 17:44:14: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
