netcdf CFS-atmos-northPacific-Vwind-2009 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:58:59 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2009/roms-cfs-atmos-Vwind-2009.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Vwind-2009.nc\n",
			"Mon Sep 10 13:44:47 2018: Time overhang added\n",
			"Mon Sep 10 13:44:43 2018: ncrcat /tmp/tp37b07c77_fec5_4000_9463_c942c05324f1.nc frc/roms-cfs-atmos-Vwind-2009.nc /tmp/tp11f34e93_4cff_4bdb_b899_3f8a56a96583.nc /tmp/tp5e583a68_802b_4bb9_a683_d96229f01396.nc\n",
			"Mon Sep 10 13:44:43 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2009.nc /tmp/tp37b07c77_fec5_4000_9463_c942c05324f1.nc\n",
			"Thu Sep  6 12:04:13 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2009_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2009.nc\n",
			"04-Oct-2017 18:10:30: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
