netcdf CFS-atmos-northPacific-lwrad-2019 {
dimensions:
	lat = 344 ;
	lon = 588 ;
	lrf_time = UNLIMITED ; // (1457 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double lrf_time(lrf_time) ;
		lrf_time:units = "day since 1900-01-01 00:00:00" ;
		lrf_time:time_origin = "01-JAN-1900 00:00:00" ;
		lrf_time:axis = "T" ;
		lrf_time:standard_name = "time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:missing_value = -1.e+34 ;
		lwrad_down:_FillValue = -1.e+34 ;
		lwrad_down:time = "lrf_time" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:long_name = "downward longwave radiation" ;
		lwrad_down:history = "From roms-cfs-atmos-lwrad-2019" ;

// global attributes:
		:history = "Mon Oct 31 12:40:29 2022: ncks -F -O -d lrf_time,2,1458 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-lwrad-2019.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-lwrad-2019.nc\n",
			"Fri Mar 27 16:04:53 2020: Time overhang added to both ends\n",
			"Fri Mar 27 16:04:44 2020: ncrcat /tmp/tpfd099217_69f6_43d2_aac4_82fafe5a1391.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-lwrad-2019.nc /tmp/tpba23c999_1bd9_460b_b0f6_709b441dde9a.nc /tmp/tp9fa7362f_4ea7_49d0_a079_26f8e7f8b800.nc\n",
			"Fri Mar 27 16:04:42 2020: ncks -F -d lrf_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-lwrad-2019.nc /tmp/tpfd099217_69f6_43d2_aac4_82fafe5a1391.nc\n",
			"FERRET V7.4   4-Mar-20" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
