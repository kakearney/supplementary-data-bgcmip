netcdf CFS-atmos-northPacific-swrad-1999 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:48:37 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1999/roms-cfs-atmos-swrad-1999.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1999/CFS-atmos-northPacific-swrad-1999.nc\n",
			"Mon Sep 10 14:03:49 2018: Time overhang added\n",
			"Mon Sep 10 14:03:48 2018: ncrcat /tmp/tpfd140b73_874a_40da_a4cf_7b49c1a71345.nc frc/roms-cfs-atmos-swrad-1999.nc /tmp/tpcb126252_3526_42b0_9372_45da67025e70.nc /tmp/tpf758ddda_f9ad_4d7c_ae39_ae2bd4e94492.nc\n",
			"Mon Sep 10 14:03:47 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-1999.nc /tmp/tpfd140b73_874a_40da_a4cf_7b49c1a71345.nc\n",
			"Thu Sep  6 10:27:28 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1999_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-1999.nc\n",
			"04-Oct-2017 17:47:59: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
