netcdf CFS-atmos-northPacific-Tair-1996 {
dimensions:
	tair_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:41:32 2022: ncks -F -O -d tair_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1996/roms-cfs-atmos-Tair-1996.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1996/CFS-atmos-northPacific-Tair-1996.nc\n",
			"Mon Sep 10 13:37:33 2018: Time overhang added\n",
			"Mon Sep 10 13:37:30 2018: ncrcat /tmp/tpfa51b3bc_64ab_486a_bc47_df10950f94a2.nc frc/roms-cfs-atmos-Tair-1996.nc /tmp/tp48e3e233_6a2d_4709_a846_6ef18cc0aab2.nc /tmp/tpffd4d4dc_7776_460a_ba96_8ec0e5653ca0.nc\n",
			"Mon Sep 10 13:37:29 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-1996.nc /tmp/tpfa51b3bc_64ab_486a_bc47_df10950f94a2.nc\n",
			"Thu Sep  6 09:57:51 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1996.nc\n",
			"Thu Sep  6 09:57:03 2018: ncks -O -F -d air_time,2,1465 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1996_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1996.nc\n",
			"04-Oct-2017 17:39:23: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
