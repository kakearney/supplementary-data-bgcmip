netcdf CFS-atmos-northPacific-Uwind-2010 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:01:45 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2010/roms-cfs-atmos-Uwind-2010.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Uwind-2010.nc\n",
			"Mon Sep 10 13:41:47 2018: Time overhang added\n",
			"Mon Sep 10 13:41:43 2018: ncrcat /tmp/tpf8354307_fee4_4b17_ba41_54ab4547ac47.nc frc/roms-cfs-atmos-Uwind-2010.nc /tmp/tp3c4da418_9836_42c5_bf93_21a53be32511.nc /tmp/tp9413ab9b_9d18_4717_86f4_341ec723d2ea.nc\n",
			"Mon Sep 10 13:41:43 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2010.nc /tmp/tpf8354307_fee4_4b17_ba41_54ab4547ac47.nc\n",
			"Thu Sep  6 12:11:01 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2010_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2010.nc\n",
			"04-Oct-2017 18:12:30: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
