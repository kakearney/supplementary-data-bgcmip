netcdf CFS-atmos-northPacific-lwrad-1999 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:47:56 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1999/roms-cfs-atmos-lwrad-1999.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1999/CFS-atmos-northPacific-lwrad-1999.nc\n",
			"Mon Sep 10 13:46:54 2018: Time overhang added\n",
			"Mon Sep 10 13:46:50 2018: ncrcat /tmp/tpa9c14284_8f92_4e4f_8076_f516d9aa139a.nc frc/roms-cfs-atmos-lwrad-1999.nc /tmp/tp8f916ea6_ffb9_4e1d_ac05_f3ea8de768c2.nc /tmp/tp4573e3ec_cc3a_4cec_8f10_ea059c2ed016.nc\n",
			"Mon Sep 10 13:46:50 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-1999.nc /tmp/tpa9c14284_8f92_4e4f_8076_f516d9aa139a.nc\n",
			"Thu Sep  6 10:26:03 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1999_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-1999.nc\n",
			"04-Oct-2017 17:47:35: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
