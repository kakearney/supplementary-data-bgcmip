netcdf CFS-atmos-northPacific-Pair-2013 {
dimensions:
	pair_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:20:35 2022: ncks -F -O -d pair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2013/roms-cfs-atmos-Pair-2013.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Pair-2013.nc\n",
			"Mon Sep 10 13:33:32 2018: Time overhang added\n",
			"Mon Sep 10 13:33:24 2018: ncrcat /tmp/tp3314662d_05a3_4840_9e40_b318dc894bc2.nc frc/roms-cfs-atmos-Pair-2013.nc /tmp/tpb5253b19_e115_4d8f_ae24_d2ea81512410.nc /tmp/tp67f6bdc4_6550_4070_83c4_6303962ddc95.nc\n",
			"Mon Sep 10 13:33:24 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2013.nc /tmp/tp3314662d_05a3_4840_9e40_b318dc894bc2.nc\n",
			"Thu Sep  6 12:51:28 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2013.nc\n",
			"Thu Sep  6 12:49:53 2018: ncks -O -F -d air_time,2,1449 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2013_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2013.nc\n",
			"04-Oct-2017 18:21:22: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
