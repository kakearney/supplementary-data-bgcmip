netcdf CFS-atmos-northPacific-Uwind-2007 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:54:09 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2007/roms-cfs-atmos-Uwind-2007.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2007/CFS-atmos-northPacific-Uwind-2007.nc\n",
			"Mon Sep 10 13:41:30 2018: Time overhang added\n",
			"Mon Sep 10 13:41:26 2018: ncrcat /tmp/tpcc45d3df_088f_4051_83ac_40ba2e6aef7b.nc frc/roms-cfs-atmos-Uwind-2007.nc /tmp/tp5d0bbf5b_5b4f_41a4_bdd6_0749f4b572c5.nc /tmp/tp2b33dfb2_7583_41c6_b10b_f03a7d57bff6.nc\n",
			"Mon Sep 10 13:41:26 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2007.nc /tmp/tpcc45d3df_088f_4051_83ac_40ba2e6aef7b.nc\n",
			"Thu Sep  6 11:47:39 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2007_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2007.nc\n",
			"04-Oct-2017 18:06:30: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
