netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2003 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:32:46 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 15:29:34 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2003/CFS-ocean-NEP-N30-bryocn-2003.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2003/CFS-ocean-ESPER-NEP-N30-brycarbon-2003.nc\n",
			"Sun Dec 25 15:15:36 2022: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad73.nc <>/final/2003/CFS-ocean-NEP-N30-bryocn-2003.nc\n",
			"Sun Dec 25 15:13:41 2022: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad01.nc\n",
			"Sun Dec 25 15:13:40 2022: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad01.nc\n",
			"Sun Dec 25 15:13:39 2022: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2003010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2003pentad01.nc\n",
			"Sun Dec 25 02:21:02 2022: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
