netcdf CFS-atmos-northPacific-rain-2020 {
dimensions:
	lat = 344 ;
	lon = 588 ;
	rain_time = UNLIMITED ; // (1447 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double rain(rain_time, lat, lon) ;
		rain:missing_value = -1.e+34 ;
		rain:_FillValue = -1.e+34 ;
		rain:time = "rain_time" ;
		rain:coordinates = "lon lat" ;
		rain:long_name = "rainfall" ;
		rain:history = "From roms-cfs-atmos-rain-2020" ;
	double rain_time(rain_time) ;
		rain_time:units = "day since 1900-01-01 00:00:00" ;
		rain_time:time_origin = "01-JAN-1900 00:00:00" ;
		rain_time:axis = "T" ;
		rain_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 13:05:21 2022: ncks -F -O -d rain_time,2,1448 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-rain-2020.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-rain-2020.nc\n",
			"Wed Jan 27 10:12:52 2021: Time overhang added to both ends\n",
			"Wed Jan 27 10:12:42 2021: ncrcat /tmp/tp13ae75da_13e8_4ba8_bc48_f2e33cd21e99.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-rain-2020.nc /tmp/tp8ece0a6d_1f1a_4f8f_98fa_fb61cd8129d1.nc /tmp/tp4134f218_f8af_4811_a94a_d77439216085.nc\n",
			"Wed Jan 27 10:12:40 2021: ncks -F -d rain_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-rain-2020.nc /tmp/tp13ae75da_13e8_4ba8_bc48_f2e33cd21e99.nc\n",
			"FERRET V7.6  26-Jan-21" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
