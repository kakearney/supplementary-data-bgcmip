netcdf CFS-atmos-northPacific-Pair-2020 {
dimensions:
	pair_time = UNLIMITED ; // (1448 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:missing_value = -1.e+34 ;
		Pair:_FillValue = -1.e+34 ;
		Pair:time = "pair_time" ;
		Pair:coordinates = "lon lat" ;
		Pair:long_name = "atmos pressure" ;
		Pair:history = "From roms-cfs-atmos-Pair-2020" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double pair_time(pair_time) ;
		pair_time:units = "day since 1900-01-01 00:00:00" ;
		pair_time:time_origin = "01-JAN-1900 00:00:00" ;
		pair_time:axis = "T" ;
		pair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:50:25 2022: ncks -F -O -d pair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Pair-2020.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Pair-2020.nc\n",
			"Wed Jan 27 10:10:36 2021: Time overhang added to both ends\n",
			"Wed Jan 27 10:10:25 2021: ncrcat /tmp/tp6a8b3833_7ae1_4753_89f0_ae8b75ac2193.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Pair-2020.nc /tmp/tp1fdc8dd6_6d37_46db_90a4_a504dde8637f.nc /tmp/tpf46f24ba_2e92_4c69_8402_89bbc8826eed.nc\n",
			"Wed Jan 27 10:10:22 2021: ncks -F -d pair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Pair-2020.nc /tmp/tp6a8b3833_7ae1_4753_89f0_ae8b75ac2193.nc\n",
			"FERRET V7.6  26-Jan-21" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
