netcdf CFS-atmos-northPacific-Uwind-2018 {
dimensions:
	wind_time = UNLIMITED ; // (1451 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:missing_value = -1.e+34 ;
		Uwind:_FillValue = -1.e+34 ;
		Uwind:time = "wind_time" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:height_above_ground1 = 10.f ;
		Uwind:long_name = "U wind" ;
		Uwind:history = "From roms-cfs-atmos-Uwind-2018" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:24:21 2022: ncks -F -O -d wind_time,2,1452 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Uwind-2018.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Uwind-2018.nc\n",
			"Thu May 30 20:49:14 2019: Time overhang added\n",
			"Thu May 30 20:49:07 2019: ncrcat /tmp/tp50ccd3b0_6546_4c54_a81a_309e59f01448.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Uwind-2018.nc /tmp/tpce974176_8ca5_4b06_a15f_99a6304a2426.nc /tmp/tp7b729133_461a_4b2a_b0e4_26078f3c1ef6.nc\n",
			"Thu May 30 20:49:07 2019: ncks -F -d wind_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Uwind-2018.nc /tmp/tp50ccd3b0_6546_4c54_a81a_309e59f01448.nc\n",
			"FERRET V7.4  29-May-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
