netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2019 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 16:52:37 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:50:01 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2019/CFS-ocean-NEP-N30-bryocn-2019.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2019/CFS-ocean-ESPER-NEP-N30-brycarbon-2019.nc\n",
			"Thu Jan 12 08:13:00 2023: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad73.nc <>/final/2019/CFS-ocean-NEP-N30-bryocn-2019.nc\n",
			"Thu Jan 12 08:08:52 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad01.nc\n",
			"Thu Jan 12 08:08:51 2023: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad01.nc\n",
			"Thu Jan 12 08:08:49 2023: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2019010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2019pentad01.nc\n",
			"Wed Jan 11 19:34:06 2023: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
