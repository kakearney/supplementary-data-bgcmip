netcdf CFS-atmos-northPacific-swrad-2009 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:59:58 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2009/roms-cfs-atmos-swrad-2009.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-swrad-2009.nc\n",
			"Mon Sep 10 14:04:11 2018: Time overhang added\n",
			"Mon Sep 10 14:04:10 2018: ncrcat /tmp/tpab075e2a_3cf5_4d0c_a47c_7e5fcd08f145.nc frc/roms-cfs-atmos-swrad-2009.nc /tmp/tpecc236e0_71d0_4b5f_93b8_0c852a08d460.nc /tmp/tp4b19fbd2_7383_487b_8a78_17132d7dfbfd.nc\n",
			"Mon Sep 10 14:04:09 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-2009.nc /tmp/tpab075e2a_3cf5_4d0c_a47c_7e5fcd08f145.nc\n",
			"Thu Sep  6 12:03:10 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2009_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-2009.nc\n",
			"04-Oct-2017 18:10:26: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
