netcdf CFS-atmos-northPacific-Tair-2010 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:00:55 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2010/roms-cfs-atmos-Tair-2010.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Tair-2010.nc\n",
			"Mon Sep 10 13:38:50 2018: Time overhang added\n",
			"Mon Sep 10 13:38:46 2018: ncrcat /tmp/tpd3f09187_6f70_4ef6_873a_321da2dec45c.nc frc/roms-cfs-atmos-Tair-2010.nc /tmp/tp572f703f_d20f_4434_9af1_22ec12c82366.nc /tmp/tp04c204f9_7b97_4470_a33c_a8d1cdc45d6a.nc\n",
			"Mon Sep 10 13:38:46 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2010.nc /tmp/tpd3f09187_6f70_4ef6_873a_321da2dec45c.nc\n",
			"Thu Sep  6 12:07:13 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2010.nc\n",
			"Thu Sep  6 12:06:17 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2010_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2010.nc\n",
			"04-Oct-2017 18:11:27: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
