netcdf CFS-atmos-northPacific-rain-2013 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	rain_time = UNLIMITED ; // (1448 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:29:47 2022: ncks -F -O -d rain_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2013/roms-cfs-atmos-rain-2013.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-rain-2013.nc\n",
			"Mon Sep 10 14:02:39 2018: Time overhang added\n",
			"Mon Sep 10 14:02:31 2018: ncrcat /tmp/tpe624bf1f_20e3_4b81_a0dd_ce4f61713896.nc frc/roms-cfs-atmos-rain-2013.nc /tmp/tp9105eaf2_dcd0_4a3a_84e6_a5a5c1e21d09.nc /tmp/tpda3dfdf6_9d54_4140_aad3_6446d2ebe779.nc\n",
			"Mon Sep 10 14:02:30 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2013.nc /tmp/tpe624bf1f_20e3_4b81_a0dd_ce4f61713896.nc\n",
			"Thu Sep  6 13:05:21 2018: ncks -O -F -d rain_time,2,1449 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2013_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2013.nc\n",
			"04-Oct-2017 18:24:34: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
