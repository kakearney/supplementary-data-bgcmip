netcdf CFS-atmos-northPacific-lwrad-1989 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	lrf_time = UNLIMITED ; // (1459 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double lrf_time(lrf_time) ;
		lrf_time:units = "day since 1900-01-01 00:00:00" ;
		lrf_time:time_origin = "01-JAN-1900 00:00:00" ;
		lrf_time:axis = "T" ;
		lrf_time:standard_name = "time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:missing_value = -1.e+34 ;
		lwrad_down:_FillValue = -1.e+34 ;
		lwrad_down:time = "lrf_time" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:long_name = "downward longwave radiation" ;
		lwrad_down:history = "From roms-cfs-atmos-lwrad-1989" ;

// global attributes:
		:history = "Fri Oct 28 16:23:56 2022: ncks -F -O -d lrf_time,2,1460 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1989/roms-cfs-atmos-lwrad-1989.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1989/CFS-atmos-northPacific-lwrad-1989.nc\n",
			"Wed Nov 20 13:55:23 2019: Time overhang added to end\n",
			"Wed Nov 20 13:55:16 2019: ncrcat /gscratch/bumblereem/bering10k/input/hindcast_cfs/1989/roms-cfs-atmos-lwrad-1989.nc /tmp/tpce4e2166_8c7e_4d20_8ef8_7ce6113c575c.nc /tmp/tp90af05d5_65a7_445e_b529_36b12252ce8b.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
