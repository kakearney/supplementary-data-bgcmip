netcdf CFS-atmos-northPacific-Tair-1995 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:37:08 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1995/roms-cfs-atmos-Tair-1995.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1995/CFS-atmos-northPacific-Tair-1995.nc\n",
			"Mon Sep 10 13:37:28 2018: Time overhang added\n",
			"Mon Sep 10 13:37:24 2018: ncrcat /tmp/tpbd848b0b_a5ef_40bc_ba04_4c393d24246f.nc frc/roms-cfs-atmos-Tair-1995.nc /tmp/tpf345f935_d6d5_4400_abd1_b0f81acd4636.nc /tmp/tp4cffbdbd_b400_492b_bd80_a9d2a980287e.nc\n",
			"Mon Sep 10 13:37:24 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-1995.nc /tmp/tpbd848b0b_a5ef_40bc_ba04_4c393d24246f.nc\n",
			"Thu Sep  6 09:50:44 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1995.nc\n",
			"Thu Sep  6 09:49:48 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1995_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1995.nc\n",
			"04-Oct-2017 17:36:52: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
