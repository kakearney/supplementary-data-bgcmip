netcdf CFS-atmos-northPacific-Vwind-2010 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:01:51 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2010/roms-cfs-atmos-Vwind-2010.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Vwind-2010.nc\n",
			"Mon Sep 10 13:44:53 2018: Time overhang added\n",
			"Mon Sep 10 13:44:49 2018: ncrcat /tmp/tpaaded371_319c_4c0a_bbef_6c922de12e44.nc frc/roms-cfs-atmos-Vwind-2010.nc /tmp/tpe2284ed7_ba64_4b8d_95f9_0439315bcd7a.nc /tmp/tpc3e750e8_589d_4775_9a95_8d304447485e.nc\n",
			"Mon Sep 10 13:44:49 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2010.nc /tmp/tpaaded371_319c_4c0a_bbef_6c922de12e44.nc\n",
			"Thu Sep  6 12:11:43 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2010_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2010.nc\n",
			"04-Oct-2017 18:12:30: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
