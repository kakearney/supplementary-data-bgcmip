netcdf CFS-atmos-northPacific-rain-2004 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1464 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:17 2022: ncks -F -O -d rain_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2004/roms-cfs-atmos-rain-2004.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2004/CFS-atmos-northPacific-rain-2004.nc\n",
			"Mon Sep 10 13:50:36 2018: Time overhang added\n",
			"Mon Sep 10 13:50:32 2018: ncrcat /tmp/tpbca762ac_4dcc_4e52_a036_c29aeb4e014c.nc frc/roms-cfs-atmos-rain-2004.nc /tmp/tpff0321e6_6132_40be_bba1_ddf757dd1bf6.nc /tmp/tp95914edf_1d5a_4a5f_aa2a_35283efe6726.nc\n",
			"Mon Sep 10 13:50:31 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2004.nc /tmp/tpbca762ac_4dcc_4e52_a036_c29aeb4e014c.nc\n",
			"Thu Sep  6 11:13:12 2018: ncks -O -F -d rain_time,2,1465 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2004_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2004.nc\n",
			"04-Oct-2017 18:01:13: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
