netcdf CFS-atmos-northPacific-Uwind-2013 {
dimensions:
	wind_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:22:52 2022: ncks -F -O -d wind_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2013/roms-cfs-atmos-Uwind-2013.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Uwind-2013.nc\n",
			"Mon Sep 10 13:42:22 2018: Time overhang added\n",
			"Mon Sep 10 13:42:13 2018: ncrcat /tmp/tp4241e0a7_629e_4171_bc8b_fe404178d742.nc frc/roms-cfs-atmos-Uwind-2013.nc /tmp/tpd51fc25a_56f5_494e_8425_ad28e28d0259.nc /tmp/tp32c1790a_628a_4f8c_9b53_b6ad3639e229.nc\n",
			"Mon Sep 10 13:42:13 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2013.nc /tmp/tp4241e0a7_629e_4171_bc8b_fe404178d742.nc\n",
			"Thu Sep  6 13:07:12 2018: ncks -O -F -d wind_time,2,1449 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2013_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2013.nc\n",
			"04-Oct-2017 18:23:31: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
