netcdf CFS-atmos-northPacific-lwrad-2001 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:50:08 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2001/roms-cfs-atmos-lwrad-2001.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2001/CFS-atmos-northPacific-lwrad-2001.nc\n",
			"Mon Sep 10 13:47:05 2018: Time overhang added\n",
			"Mon Sep 10 13:47:01 2018: ncrcat /tmp/tp628ce620_2275_4842_bbee_4a1453d58a14.nc frc/roms-cfs-atmos-lwrad-2001.nc /tmp/tp9e22a8ca_2eb6_4800_a709_569a3cb94e09.nc /tmp/tp3f614914_5e38_42da_838d_6b8ac25a885b.nc\n",
			"Mon Sep 10 13:47:01 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2001.nc /tmp/tp628ce620_2275_4842_bbee_4a1453d58a14.nc\n",
			"Thu Sep  6 10:44:29 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2001_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2001.nc\n",
			"04-Oct-2017 17:52:45: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
