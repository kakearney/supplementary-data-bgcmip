netcdf CFS-atmos-northPacific-Vwind-2002 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:28 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2002/roms-cfs-atmos-Vwind-2002.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2002/CFS-atmos-northPacific-Vwind-2002.nc\n",
			"Mon Sep 10 13:44:07 2018: Time overhang added\n",
			"Mon Sep 10 13:44:03 2018: ncrcat /tmp/tp853e9d54_f6fe_4cfd_b455_855b2bd93936.nc frc/roms-cfs-atmos-Vwind-2002.nc /tmp/tp478dbbb7_cadf_42f4_a133_75e43977e989.nc /tmp/tp88208067_8e1c_4698_9cba_955d93ede110.nc\n",
			"Mon Sep 10 13:44:03 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2002.nc /tmp/tp853e9d54_f6fe_4cfd_b455_855b2bd93936.nc\n",
			"Thu Sep  6 10:57:53 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2002_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2002.nc\n",
			"04-Oct-2017 17:56:02: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
