netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-1991 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 14:28:01 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 14:26:21 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1991/CFS-ocean-Bering10K-N30-bryocn-1991.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1991/CFS-ocean-ESPER-Bering10K-N30-brycarbon-1991.nc\n",
			"Tue Dec 13 06:22:28 2022: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad73.nc <>/final/1991/CFS-ocean-Bering10K-N30-bryocn-1991.nc\n",
			"Tue Dec 13 06:21:44 2022: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad01.nc\n",
			"Tue Dec 13 06:21:44 2022: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1991010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1991pentad01.nc\n",
			"Mon Dec 12 10:30:29 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
