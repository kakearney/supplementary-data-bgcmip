netcdf CFS-atmos-northPacific-Qair-2019 {
dimensions:
	qair_time = UNLIMITED ; // (1457 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:missing_value = -1.e+34 ;
		Qair:_FillValue = -1.e+34 ;
		Qair:time = "qair_time" ;
		Qair:coordinates = "lon lat" ;
		Qair:height_above_ground = 2.f ;
		Qair:long_name = "specific humidity" ;
		Qair:history = "From roms-cfs-atmos-Qair-2019" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double qair_time(qair_time) ;
		qair_time:units = "day since 1900-01-01 00:00:00" ;
		qair_time:time_origin = "01-JAN-1900 00:00:00" ;
		qair_time:axis = "T" ;
		qair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:36:52 2022: ncks -F -O -d qair_time,2,1458 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Qair-2019.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Qair-2019.nc\n",
			"Fri Mar 27 16:03:34 2020: Time overhang added to both ends\n",
			"Fri Mar 27 16:03:25 2020: ncrcat /tmp/tp7327cf5a_e2b0_4295_9712_213d5512df26.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Qair-2019.nc /tmp/tp9b7550fd_ac5a_4b25_875e_49b4b7db0b79.nc /tmp/tp96847b6a_a282_4c90_a2b5_c89304757f05.nc\n",
			"Fri Mar 27 16:03:24 2020: ncks -F -d qair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Qair-2019.nc /tmp/tp7327cf5a_e2b0_4295_9712_213d5512df26.nc\n",
			"FERRET V7.4   4-Mar-20" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
