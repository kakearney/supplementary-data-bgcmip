netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-2022 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 17:04:40 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 17:03:04 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2022/CFS-ocean-Bering10K-N30-bryocn-2022.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2022/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2022.nc\n",
			"Sun Jan 15 19:13:25 2023: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad73.nc <>/final/2022/CFS-ocean-Bering10K-N30-bryocn-2022.nc\n",
			"Sun Jan 15 19:11:51 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad01.nc\n",
			"Sun Jan 15 19:11:51 2023: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad01.nc\n",
			"Sun Jan 15 19:11:51 2023: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2022010512.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2022pentad01.nc\n",
			"Fri Jan 13 10:38:07 2023: CFS data added\n",
			"Tue Dec 20 15:09:11 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
