netcdf CFS-atmos-northPacific-Qair-2020 {
dimensions:
	qair_time = UNLIMITED ; // (1448 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:missing_value = -1.e+34 ;
		Qair:_FillValue = -1.e+34 ;
		Qair:time = "qair_time" ;
		Qair:coordinates = "lon lat" ;
		Qair:height_above_ground = 2.f ;
		Qair:long_name = "specific humidity" ;
		Qair:history = "From roms-cfs-atmos-Qair-2020" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double qair_time(qair_time) ;
		qair_time:units = "day since 1900-01-01 00:00:00" ;
		qair_time:time_origin = "01-JAN-1900 00:00:00" ;
		qair_time:axis = "T" ;
		qair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:51:22 2022: ncks -F -O -d qair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Qair-2020.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Qair-2020.nc\n",
			"Wed Jan 27 10:10:59 2021: Time overhang added to both ends\n",
			"Wed Jan 27 10:10:49 2021: ncrcat /tmp/tpe12aab1c_0ba4_428d_b78f_8ace4510ef78.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Qair-2020.nc /tmp/tp9f4444ef_3a60_4c01_bc38_6b598998db8a.nc /tmp/tpc989bf29_47af_44bb_9760_30144abb1e89.nc\n",
			"Wed Jan 27 10:10:48 2021: ncks -F -d qair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Qair-2020.nc /tmp/tpe12aab1c_0ba4_428d_b78f_8ace4510ef78.nc\n",
			"FERRET V7.6  26-Jan-21" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
