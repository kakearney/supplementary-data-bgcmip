netcdf CFS-atmos-northPacific-Uwind-1996 {
dimensions:
	wind_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:41:38 2022: ncks -F -O -d wind_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1996/roms-cfs-atmos-Uwind-1996.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1996/CFS-atmos-northPacific-Uwind-1996.nc\n",
			"Mon Sep 10 13:40:29 2018: Time overhang added\n",
			"Mon Sep 10 13:40:26 2018: ncrcat /tmp/tp9a092c92_d800_4ce6_a452_158db4fd64ac.nc frc/roms-cfs-atmos-Uwind-1996.nc /tmp/tpd8b3657f_3f9d_4ab4_988f_3de858b62490.nc /tmp/tpb0b5843d_2900_4347_a483_1b143bdd61f2.nc\n",
			"Mon Sep 10 13:40:25 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-1996.nc /tmp/tp9a092c92_d800_4ce6_a452_158db4fd64ac.nc\n",
			"Thu Sep  6 10:01:28 2018: ncks -O -F -d wind_time,2,1465 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1996_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-1996.nc\n",
			"04-Oct-2017 17:40:44: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
