netcdf CFS-atmos-northPacific-Qair-2005 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:33 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2005/roms-cfs-atmos-Qair-2005.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2005/CFS-atmos-northPacific-Qair-2005.nc\n",
			"Mon Sep 10 13:35:27 2018: Time overhang added\n",
			"Mon Sep 10 13:35:24 2018: ncrcat /tmp/tp0f8721db_0265_466c_9208_ec74ebaf0784.nc frc/roms-cfs-atmos-Qair-2005.nc /tmp/tp52dcd03f_3570_4a2b_99ea_005c03fa8d50.nc /tmp/tp96c18165_258c_416b_af70_0a5cdf9fadc9.nc\n",
			"Mon Sep 10 13:35:23 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2005.nc /tmp/tp0f8721db_0265_466c_9208_ec74ebaf0784.nc\n",
			"Thu Sep  6 11:20:42 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2005.nc\n",
			"Thu Sep  6 11:19:44 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2005_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2005.nc\n",
			"04-Oct-2017 18:01:29: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
