netcdf CFS-atmos-northPacific-rain-1995 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:40:28 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1995/roms-cfs-atmos-rain-1995.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1995/CFS-atmos-northPacific-rain-1995.nc\n",
			"Mon Sep 10 13:49:43 2018: Time overhang added\n",
			"Mon Sep 10 13:49:40 2018: ncrcat /tmp/tpda14aac6_c27c_4290_a6b0_4b972c1b28af.nc frc/roms-cfs-atmos-rain-1995.nc /tmp/tpd940059c_326e_4857_a227_6317e4a00b83.nc /tmp/tp5b754a01_67d4_4541_b170_629e01b8a7ce.nc\n",
			"Mon Sep 10 13:49:39 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-1995.nc /tmp/tpda14aac6_c27c_4290_a6b0_4b972c1b28af.nc\n",
			"Thu Sep  6 09:53:22 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1995_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-1995.nc\n",
			"04-Oct-2017 17:39:00: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
