netcdf CFS-atmos-northPacific-lwrad-1984 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double lrf_time(lrf_time) ;
		lrf_time:units = "day since 1900-01-01 00:00:00" ;
		lrf_time:time_origin = "01-JAN-1900 00:00:00" ;
		lrf_time:axis = "T" ;
		lrf_time:standard_name = "time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:missing_value = -1.e+34 ;
		lwrad_down:_FillValue = -1.e+34 ;
		lwrad_down:time = "lrf_time" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:long_name = "downward longwave radiation" ;
		lwrad_down:history = "From roms-cfs-atmos-lwrad-1984" ;

// global attributes:
		:history = "Thu Nov  3 15:35:06 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-lwrad-1984.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1984/CFS-atmos-northPacific-lwrad-1984.nc\n",
			"Wed Nov 20 13:45:00 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:44:56 2019: ncrcat /tmp/tp2dba0511_e9fb_43dc_9178_5abf7688c332.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-lwrad-1984.nc /tmp/tp9ae47eec_169c_498c_a933_f8f73e157fd6.nc /tmp/tp70febce4_97cb_4f82_8fcb_63d4b6fce644.nc\n",
			"Wed Nov 20 13:44:54 2019: ncks -F -d lrf_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-lwrad-1984.nc /tmp/tp2dba0511_e9fb_43dc_9178_5abf7688c332.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
