netcdf CFS-atmos-northPacific-lwrad-2004 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1464 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:08 2022: ncks -F -O -d lrf_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2004/roms-cfs-atmos-lwrad-2004.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2004/CFS-atmos-northPacific-lwrad-2004.nc\n",
			"Mon Sep 10 13:47:22 2018: Time overhang added\n",
			"Mon Sep 10 13:47:18 2018: ncrcat /tmp/tp6d6b5ad4_eced_4d6d_aba2_0121390c8b2b.nc frc/roms-cfs-atmos-lwrad-2004.nc /tmp/tp8307304d_37b4_47a9_b37f_6ba3c294f0a6.nc /tmp/tp06c9e8d5_cc7e_4d40_a292_6d8257fe7872.nc\n",
			"Mon Sep 10 13:47:18 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2004.nc /tmp/tp6d6b5ad4_eced_4d6d_aba2_0121390c8b2b.nc\n",
			"Thu Sep  6 11:12:26 2018: ncks -O -F -d lrf_time,2,1465 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2004_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2004.nc\n",
			"04-Oct-2017 18:00:17: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
