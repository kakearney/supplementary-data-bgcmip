netcdf CFS-atmos-northPacific-Vwind-2007 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:54:20 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2007/roms-cfs-atmos-Vwind-2007.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2007/CFS-atmos-northPacific-Vwind-2007.nc\n",
			"Mon Sep 10 13:44:36 2018: Time overhang added\n",
			"Mon Sep 10 13:44:32 2018: ncrcat /tmp/tp7c3f75a8_81cf_4a98_b03c_697d4cbd9b1a.nc frc/roms-cfs-atmos-Vwind-2007.nc /tmp/tp5402b4a6_2662_4843_a4e6_444356bad2dc.nc /tmp/tp8f421545_1886_49a8_8427_73c0421276b1.nc\n",
			"Mon Sep 10 13:44:31 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2007.nc /tmp/tp7c3f75a8_81cf_4a98_b03c_697d4cbd9b1a.nc\n",
			"Thu Sep  6 11:48:40 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2007_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2007.nc\n",
			"04-Oct-2017 18:06:30: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
