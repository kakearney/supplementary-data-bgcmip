netcdf CFS-atmos-northPacific-rain-2005 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:52:08 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2005/roms-cfs-atmos-rain-2005.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2005/CFS-atmos-northPacific-rain-2005.nc\n",
			"Mon Sep 10 13:50:47 2018: Time overhang added\n",
			"Mon Sep 10 13:50:43 2018: ncrcat /tmp/tp911ec755_a904_4161_993a_87f7a731ab18.nc frc/roms-cfs-atmos-rain-2005.nc /tmp/tpd0e6e40d_4c01_4c49_bc0a_13474be005e9.nc /tmp/tpd630a812_3026_4ff3_a607_2c215a7fc0a5.nc\n",
			"Mon Sep 10 13:50:42 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2005.nc /tmp/tp911ec755_a904_4161_993a_87f7a731ab18.nc\n",
			"Thu Sep  6 11:22:28 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2005_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2005.nc\n",
			"04-Oct-2017 18:03:10: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
