netcdf CFS-atmos-northPacific-Pair-2016 {
dimensions:
	pair_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Mon Oct 31 11:53:19 2022: ncks -F -O -d pair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2016/roms-cfs-atmos-Pair-2016.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Pair-2016.nc\n",
			"Mon Sep 10 13:34:06 2018: Time overhang added\n",
			"Mon Sep 10 13:33:58 2018: ncrcat /tmp/tp67c7de34_1100_400e_8678_4484b35d58e1.nc frc/roms-cfs-atmos-Pair-2016.nc /tmp/tp00b85720_98be_4205_87af_c1269631ca6e.nc /tmp/tpafd88ea4_28c7_4f34_973a_de30a20143c3.nc\n",
			"Mon Sep 10 13:33:57 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2016.nc /tmp/tp67c7de34_1100_400e_8678_4484b35d58e1.nc\n",
			"Thu Sep  6 13:59:35 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2016.nc\n",
			"Thu Sep  6 13:57:31 2018: ncks -O -F -d air_time,2,1449 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2016_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2016.nc\n",
			"04-Oct-2017 18:32:42: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
