netcdf CFS-atmos-northPacific-rain-2008 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1464 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:57:39 2022: ncks -F -O -d rain_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2008/roms-cfs-atmos-rain-2008.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2008/CFS-atmos-northPacific-rain-2008.nc\n",
			"Mon Sep 10 13:51:04 2018: Time overhang added\n",
			"Mon Sep 10 13:51:01 2018: ncrcat /tmp/tpb230f202_2b9a_43bd_91d0_9b865ad8b05a.nc frc/roms-cfs-atmos-rain-2008.nc /tmp/tpbf463a7a_e8d1_4886_b142_0f06796011a7.nc /tmp/tp38ba239c_624a_4554_a0a1_a8f65bfe0325.nc\n",
			"Mon Sep 10 13:51:00 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2008.nc /tmp/tpb230f202_2b9a_43bd_91d0_9b865ad8b05a.nc\n",
			"Thu Sep  6 11:54:56 2018: ncks -O -F -d rain_time,2,1465 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2008_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2008.nc\n",
			"04-Oct-2017 18:09:08: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
