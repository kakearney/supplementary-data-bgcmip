netcdf CFS-atmos-northPacific-Tair-2019 {
dimensions:
	tair_time = UNLIMITED ; // (1457 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:missing_value = -1.e+34 ;
		Tair:_FillValue = -1.e+34 ;
		Tair:time = "tair_time" ;
		Tair:coordinates = "lon lat" ;
		Tair:height_above_ground = 2.f ;
		Tair:long_name = "surface air temperature" ;
		Tair:history = "From roms-cfs-atmos-Tair-2019" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double tair_time(tair_time) ;
		tair_time:units = "day since 1900-01-01 00:00:00" ;
		tair_time:time_origin = "01-JAN-1900 00:00:00" ;
		tair_time:axis = "T" ;
		tair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:37:46 2022: ncks -F -O -d tair_time,2,1458 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Tair-2019.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Tair-2019.nc\n",
			"Fri Mar 27 16:03:55 2020: Time overhang added to both ends\n",
			"Fri Mar 27 16:03:44 2020: ncrcat /tmp/tpd13120fd_71a4_45a3_a9f3_7622015ed848.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Tair-2019.nc /tmp/tp74e7052e_d94e_4242_8daa_4edf67175489.nc /tmp/tpec03cc57_9ed8_4a7e_8ce7_b791ac56f86b.nc\n",
			"Fri Mar 27 16:03:42 2020: ncks -F -d tair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Tair-2019.nc /tmp/tpd13120fd_71a4_45a3_a9f3_7622015ed848.nc\n",
			"FERRET V7.4   4-Mar-20" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
