netcdf CFS-atmos-northPacific-Uwind-2001 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:49:54 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2001/roms-cfs-atmos-Uwind-2001.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2001/CFS-atmos-northPacific-Uwind-2001.nc\n",
			"Mon Sep 10 13:40:57 2018: Time overhang added\n",
			"Mon Sep 10 13:40:53 2018: ncrcat /tmp/tpc0867f42_1453_449b_8a5b_8f6d0c66b720.nc frc/roms-cfs-atmos-Uwind-2001.nc /tmp/tp1652bb34_9aad_44f9_8f12_0f6ab6b12326.nc /tmp/tp85200d67_2f22_4942_aa10_e98ea7a5e6f8.nc\n",
			"Mon Sep 10 13:40:53 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2001.nc /tmp/tpc0867f42_1453_449b_8a5b_8f6d0c66b720.nc\n",
			"Thu Sep  6 10:46:50 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2001_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2001.nc\n",
			"04-Oct-2017 17:53:12: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
