netcdf CFS-atmos-northPacific-Pair-2021 {
dimensions:
	pair_time = UNLIMITED ; // (1431 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:missing_value = -1.e+34 ;
		Pair:_FillValue = -1.e+34 ;
		Pair:time = "pair_time" ;
		Pair:coordinates = "lon lat" ;
		Pair:long_name = "atmos pressure" ;
		Pair:history = "From roms-cfs-atmos-Pair-2021" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double pair_time(pair_time) ;
		pair_time:units = "day since 1900-01-01 00:00:00" ;
		pair_time:time_origin = "01-JAN-1900 00:00:00" ;
		pair_time:axis = "T" ;
		pair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 13:06:28 2022: ncks -F -O -d pair_time,2,1432 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2021/roms-cfs-atmos-Pair-2021.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2021/CFS-atmos-northPacific-Pair-2021.nc\n",
			"Fri May 06 13:50:26 2022: Time overhang added to end\n",
			"Fri May  6 13:50:15 2022: ncrcat /gscratch/bumblereem/bering10k/input/hindcast_cfs/2021/roms-cfs-atmos-Pair-2021.nc /tmp/tp6e680bb5_1335_4ab2_83c5_93e899d03df5.nc /tmp/tpb17c921c_2397_4773_bdf9_c04f5a2c2b01.nc\n",
			"FERRET V7.6  20-Jan-22" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
