netcdf CFS-atmos-northPacific-lwrad-1986 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double lrf_time(lrf_time) ;
		lrf_time:units = "day since 1900-01-01 00:00:00" ;
		lrf_time:time_origin = "01-JAN-1900 00:00:00" ;
		lrf_time:axis = "T" ;
		lrf_time:standard_name = "time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:missing_value = -1.e+34 ;
		lwrad_down:_FillValue = -1.e+34 ;
		lwrad_down:time = "lrf_time" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:long_name = "downward longwave radiation" ;
		lwrad_down:history = "From roms-cfs-atmos-lwrad-1986" ;

// global attributes:
		:history = "Fri Oct 28 16:19:57 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-lwrad-1986.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1986/CFS-atmos-northPacific-lwrad-1986.nc\n",
			"Wed Nov 20 13:49:00 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:48:54 2019: ncrcat /tmp/tpf3d61425_db5f_444d_af0c_8ce8d80ab155.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-lwrad-1986.nc /tmp/tp8e6ff3ff_005b_4d24_904f_1b138b734434.nc /tmp/tp37725255_9cdd_48d5_b9c1_224a1de7d60c.nc\n",
			"Wed Nov 20 13:48:52 2019: ncks -F -d lrf_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-lwrad-1986.nc /tmp/tpf3d61425_db5f_444d_af0c_8ce8d80ab155.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
