netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-2013 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 16:20:23 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:18:48 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2013/CFS-ocean-Bering10K-N30-bryocn-2013.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2013/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2013.nc\n",
			"Sun Jan  8 19:52:00 2023: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad73.nc <>/final/2013/CFS-ocean-Bering10K-N30-bryocn-2013.nc\n",
			"Sun Jan  8 19:50:50 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad01.nc\n",
			"Sun Jan  8 19:50:50 2023: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad01.nc\n",
			"Sun Jan  8 19:50:49 2023: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2013010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2013pentad01.nc\n",
			"Sun Jan 08 06:23:27 2023: CFS data added\n",
			"Tue Dec 20 15:09:11 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
