netcdf CFS-atmos-northPacific-swrad-1995 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:41:15 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1995/roms-cfs-atmos-swrad-1995.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1995/CFS-atmos-northPacific-swrad-1995.nc\n",
			"Mon Sep 10 14:03:40 2018: Time overhang added\n",
			"Mon Sep 10 14:03:39 2018: ncrcat /tmp/tp9ec04c63_bd48_4c08_b7a9_6f188fc99850.nc frc/roms-cfs-atmos-swrad-1995.nc /tmp/tp1d2e5cbb_a933_4e98_b430_41fdcb3bbb49.nc /tmp/tp03c5caba_d53c_4fb5_b498_f8e205b2d934.nc\n",
			"Mon Sep 10 14:03:39 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-1995.nc /tmp/tp9ec04c63_bd48_4c08_b7a9_6f188fc99850.nc\n",
			"Thu Sep  6 09:53:56 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1995_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-1995.nc\n",
			"04-Oct-2017 17:38:12: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
