netcdf CFS-atmos-northPacific-rain-2019 {
dimensions:
	lat = 344 ;
	lon = 588 ;
	rain_time = UNLIMITED ; // (1457 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double rain(rain_time, lat, lon) ;
		rain:missing_value = -1.e+34 ;
		rain:_FillValue = -1.e+34 ;
		rain:time = "rain_time" ;
		rain:coordinates = "lon lat" ;
		rain:long_name = "rainfall" ;
		rain:history = "From roms-cfs-atmos-rain-2019" ;
	double rain_time(rain_time) ;
		rain_time:units = "day since 1900-01-01 00:00:00" ;
		rain_time:time_origin = "01-JAN-1900 00:00:00" ;
		rain_time:axis = "T" ;
		rain_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:49:28 2022: ncks -F -O -d rain_time,2,1458 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-rain-2019.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-rain-2019.nc\n",
			"Fri Mar 27 16:05:30 2020: Time overhang added to both ends\n",
			"Fri Mar 27 16:05:21 2020: ncrcat /tmp/tpc972c67e_f397_44e9_acbc_f3d2ab1d1a5e.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-rain-2019.nc /tmp/tpe7cd279f_3f89_4f80_a25b_6787b9b2b4ef.nc /tmp/tpb5825d10_b8d9_4e2e_9f7d_31aa5e43dc4a.nc\n",
			"Fri Mar 27 16:05:19 2020: ncks -F -d rain_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-rain-2019.nc /tmp/tpc972c67e_f397_44e9_acbc_f3d2ab1d1a5e.nc\n",
			"FERRET V7.4   4-Mar-20" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
