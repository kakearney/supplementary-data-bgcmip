netcdf CFS-atmos-northPacific-Tair-2011 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:03:48 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2011/roms-cfs-atmos-Tair-2011.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Tair-2011.nc\n",
			"Thu Sep 13 10:47:58 2018: Time overhang added\n",
			"Thu Sep 13 10:47:51 2018: ncrcat /tmp/tpe47609c7_b3a2_4a65_ac5d_ecf46edb6c8f.nc frc/roms-cfs-atmos-Tair-2011.nc /tmp/tp4f831a62_34a7_4a5f_b161_13f4c3f1837a.nc /tmp/tp25a4f09d_9076_4977_9428_44629aa00eaa.nc\n",
			"Thu Sep 13 10:47:51 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2011.nc /tmp/tpe47609c7_b3a2_4a65_ac5d_ecf46edb6c8f.nc\n",
			"Thu Sep 13 10:41:32 2018: ncrename -d air_time,tair_time -v air_time,tair_time ./frc/roms-cfs-atmos-Tair-2011.nc\n",
			"Thu Sep 13 10:41:22 2018: ncks -O -F -d air_time,2,1461 -v Tair ./frc/Old/corecfs_2011_air.nc ./frc/roms-cfs-atmos-Tair-2011.nc\n",
			"04-Oct-2017 18:13:26: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
