netcdf CFS-atmos-northPacific-Pair-2008 {
dimensions:
	pair_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:55:08 2022: ncks -F -O -d pair_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2008/roms-cfs-atmos-Pair-2008.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2008/CFS-atmos-northPacific-Pair-2008.nc\n",
			"Mon Sep 10 13:32:49 2018: Time overhang added\n",
			"Mon Sep 10 13:32:46 2018: ncrcat /tmp/tpa08b9479_43e2_4143_b32d_2a198e562446.nc frc/roms-cfs-atmos-Pair-2008.nc /tmp/tpd9e4d5c1_91ff_4ec6_a869_b68b841b2e6e.nc /tmp/tp90aa37d9_1614_41b6_922e_8685663ed986.nc\n",
			"Mon Sep 10 13:32:45 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2008.nc /tmp/tpa08b9479_43e2_4143_b32d_2a198e562446.nc\n",
			"Thu Sep  6 11:50:49 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2008.nc\n",
			"Thu Sep  6 11:49:46 2018: ncks -O -F -d air_time,2,1465 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2008_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2008.nc\n",
			"04-Oct-2017 18:07:27: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
