netcdf CFS-atmos-northPacific-Pair-1998 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:49 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1998/roms-cfs-atmos-Pair-1998.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1998/CFS-atmos-northPacific-Pair-1998.nc\n",
			"Mon Sep 10 13:31:54 2018: Time overhang added\n",
			"Mon Sep 10 13:31:50 2018: ncrcat /tmp/tp42e75023_f150_44b4_ab9b_f6f0a5c10542.nc frc/roms-cfs-atmos-Pair-1998.nc /tmp/tp3a6d90bb_dc79_4444_9748_ce89b9cfb343.nc /tmp/tpa5647a01_f969_4823_9567_2f36ba15f130.nc\n",
			"Mon Sep 10 13:31:48 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-1998.nc /tmp/tp42e75023_f150_44b4_ab9b_f6f0a5c10542.nc\n",
			"Thu Sep  6 10:13:57 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1998.nc\n",
			"Thu Sep  6 10:13:00 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1998_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1998.nc\n",
			"04-Oct-2017 17:44:14: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
