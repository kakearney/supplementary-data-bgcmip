netcdf CFS-atmos-northPacific-lwrad-1988 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double lrf_time(lrf_time) ;
		lrf_time:units = "day since 1900-01-01 00:00:00" ;
		lrf_time:time_origin = "01-JAN-1900 00:00:00" ;
		lrf_time:axis = "T" ;
		lrf_time:standard_name = "time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:missing_value = -1.e+34 ;
		lwrad_down:_FillValue = -1.e+34 ;
		lwrad_down:time = "lrf_time" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:long_name = "downward longwave radiation" ;
		lwrad_down:history = "From roms-cfs-atmos-lwrad-1988" ;

// global attributes:
		:history = "Fri Oct 28 16:21:39 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1988/roms-cfs-atmos-lwrad-1988.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1988/CFS-atmos-northPacific-lwrad-1988.nc\n",
			"Wed Nov 20 13:53:19 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:53:14 2019: ncrcat /tmp/tp25b5061d_0237_4d88_9401_d7619d29459e.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1988/roms-cfs-atmos-lwrad-1988.nc /tmp/tpe9ca0743_3bfd_4865_97f0_145776a2daaf.nc /tmp/tp2f368597_a526_4653_bcf5_f5ed3ef1a02e.nc\n",
			"Wed Nov 20 13:53:12 2019: ncks -F -d lrf_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1988/roms-cfs-atmos-lwrad-1988.nc /tmp/tp25b5061d_0237_4d88_9401_d7619d29459e.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
