netcdf CFS-atmos-northPacific-rain-1992 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double rain(rain_time, lat, lon) ;
		rain:missing_value = -1.e+34 ;
		rain:_FillValue = -1.e+34 ;
		rain:time = "rain_time" ;
		rain:coordinates = "lon lat" ;
		rain:long_name = "rainfall" ;
		rain:history = "From roms-cfs-atmos-rain-1992" ;
	double rain_time(rain_time) ;
		rain_time:units = "day since 1900-01-01 00:00:00" ;
		rain_time:time_origin = "01-JAN-1900 00:00:00" ;
		rain_time:axis = "T" ;
		rain_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:30:59 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1992/roms-cfs-atmos-rain-1992.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1992/CFS-atmos-northPacific-rain-1992.nc\n",
			"Wed Nov 20 14:02:02 2019: Time overhang added to both ends\n",
			"Wed Nov 20 14:01:58 2019: ncrcat /tmp/tp83aa9cf0_5466_4eac_a99e_ea1ffaf50748.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1992/roms-cfs-atmos-rain-1992.nc /tmp/tp59eb9b1a_57fa_462f_a6e3_4aa936941336.nc /tmp/tp93c90653_1609_4b7c_89d6_49da60ebebb2.nc\n",
			"Wed Nov 20 14:01:56 2019: ncks -F -d rain_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1992/roms-cfs-atmos-rain-1992.nc /tmp/tp83aa9cf0_5466_4eac_a99e_ea1ffaf50748.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
