netcdf CFS-atmos-northPacific-Qair-1999 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:47:27 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1999/roms-cfs-atmos-Qair-1999.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1999/CFS-atmos-northPacific-Qair-1999.nc\n",
			"Mon Sep 10 13:34:55 2018: Time overhang added\n",
			"Mon Sep 10 13:34:51 2018: ncrcat /tmp/tp86030d0f_af81_42b3_a86f_28d47066afb6.nc frc/roms-cfs-atmos-Qair-1999.nc /tmp/tp193aaefe_25f8_41b2_8f03_dfb97e1ff073.nc /tmp/tp86e2944c_6b0b_4d97_bedd_17fb8f897bb2.nc\n",
			"Mon Sep 10 13:34:51 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-1999.nc /tmp/tp86030d0f_af81_42b3_a86f_28d47066afb6.nc\n",
			"Thu Sep  6 10:25:14 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-1999.nc\n",
			"Thu Sep  6 10:24:23 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1999_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-1999.nc\n",
			"04-Oct-2017 17:46:41: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
