netcdf CFS-atmos-northPacific-Vwind-2012 {
dimensions:
	wind_time = UNLIMITED ; // (1464 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:15:00 2022: ncks -F -O -d wind_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2012/roms-cfs-atmos-Vwind-2012.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Vwind-2012.nc\n",
			"Mon Sep 10 13:45:15 2018: Time overhang added\n",
			"Mon Sep 10 13:45:07 2018: ncrcat /tmp/tp4e6acd16_3ba1_4fee_bad7_c54615cab8d2.nc frc/roms-cfs-atmos-Vwind-2012.nc /tmp/tpb05bcc4e_1dc8_493c_8d90_6100b8a02a92.nc /tmp/tpf1ebe4c8_99ce_48e8_a2c0_c45ffda5ede1.nc\n",
			"Mon Sep 10 13:45:06 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2012.nc /tmp/tp4e6acd16_3ba1_4fee_bad7_c54615cab8d2.nc\n",
			"Thu Sep  6 12:48:10 2018: ncks -O -F -d wind_time,2,1465 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2012_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2012.nc\n",
			"04-Oct-2017 18:19:43: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
