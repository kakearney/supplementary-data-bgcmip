netcdf CFS-atmos-northPacific-Vwind-2004 {
dimensions:
	wind_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:00 2022: ncks -F -O -d wind_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2004/roms-cfs-atmos-Vwind-2004.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2004/CFS-atmos-northPacific-Vwind-2004.nc\n",
			"Mon Sep 10 13:44:18 2018: Time overhang added\n",
			"Mon Sep 10 13:44:15 2018: ncrcat /tmp/tp2bf7e72b_a98a_4863_acdb_000dcda6d3e7.nc frc/roms-cfs-atmos-Vwind-2004.nc /tmp/tpf00e7cfe_fd38_4aee_887e_cf07320da452.nc /tmp/tp1eb45189_0b2b_4a0c_b058_e57c5d10f15f.nc\n",
			"Mon Sep 10 13:44:14 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2004.nc /tmp/tp2bf7e72b_a98a_4863_acdb_000dcda6d3e7.nc\n",
			"Thu Sep  6 11:15:15 2018: ncks -O -F -d wind_time,2,1465 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2004_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2004.nc\n",
			"04-Oct-2017 18:00:38: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
