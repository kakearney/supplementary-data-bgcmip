netcdf CFS-atmos-northPacific-swrad-2003 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:17:38 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2003/roms-cfs-atmos-swrad-2003.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2003/CFS-atmos-northPacific-swrad-2003.nc\n",
			"Mon Sep 10 14:03:57 2018: Time overhang added\n",
			"Mon Sep 10 14:03:56 2018: ncrcat /tmp/tp4d26a383_7efe_45ad_b5a3_1eb4b02bd24b.nc frc/roms-cfs-atmos-swrad-2003.nc /tmp/tpca2dc51a_4bda_44bd_b735_2390a0514d76.nc /tmp/tp876c5da8_ffdf_4c90_9bbe_6b7fec253540.nc\n",
			"Mon Sep 10 14:03:55 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-2003.nc /tmp/tp4d26a383_7efe_45ad_b5a3_1eb4b02bd24b.nc\n",
			"Thu Sep  6 11:05:37 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2003_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-2003.nc\n",
			"04-Oct-2017 17:58:21: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
