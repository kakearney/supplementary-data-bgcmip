netcdf CFS-atmos-northPacific-Uwind-2008 {
dimensions:
	wind_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:56:35 2022: ncks -F -O -d wind_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2008/roms-cfs-atmos-Uwind-2008.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2008/CFS-atmos-northPacific-Uwind-2008.nc\n",
			"Mon Sep 10 13:41:36 2018: Time overhang added\n",
			"Mon Sep 10 13:41:32 2018: ncrcat /tmp/tpf439f9b4_941c_4f48_aa10_5d84849699d8.nc frc/roms-cfs-atmos-Uwind-2008.nc /tmp/tp35f7564e_0f04_4523_8f31_82e4a95bfbae.nc /tmp/tpa21d6914_28cb_4055_9bc4_f9eed750a9d3.nc\n",
			"Mon Sep 10 13:41:32 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2008.nc /tmp/tpf439f9b4_941c_4f48_aa10_5d84849699d8.nc\n",
			"Thu Sep  6 11:55:54 2018: ncks -O -F -d wind_time,2,1465 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2008_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2008.nc\n",
			"04-Oct-2017 18:08:30: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
