netcdf CFS-atmos-northPacific-lwrad-2012 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	lrf_time = UNLIMITED ; // (1464 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:15:13 2022: ncks -F -O -d lrf_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2012/roms-cfs-atmos-lwrad-2012.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-lwrad-2012.nc\n",
			"Mon Sep 10 13:48:19 2018: Time overhang added\n",
			"Mon Sep 10 13:48:10 2018: ncrcat /tmp/tpd5885873_0afa_4fd7_8f52_777ed91b7abd.nc frc/roms-cfs-atmos-lwrad-2012.nc /tmp/tpd485d71d_eb9c_46db_9d33_6a2d1cf2aff6.nc /tmp/tpd71ec609_fddb_400f_9588_d42807ecd4f9.nc\n",
			"Mon Sep 10 13:48:10 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2012.nc /tmp/tpd5885873_0afa_4fd7_8f52_777ed91b7abd.nc\n",
			"Thu Sep  6 12:43:40 2018: ncks -O -F -d lrf_time,2,1465 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2012_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2012.nc\n",
			"04-Oct-2017 18:18:52: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
