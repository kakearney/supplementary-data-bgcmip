netcdf CFS-atmos-northPacific-Pair-2001 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:49:33 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2001/roms-cfs-atmos-Pair-2001.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2001/CFS-atmos-northPacific-Pair-2001.nc\n",
			"Mon Sep 10 13:32:12 2018: Time overhang added\n",
			"Mon Sep 10 13:32:09 2018: ncrcat /tmp/tpf43628e7_83d0_4a16_bd5a_42915d7abb03.nc frc/roms-cfs-atmos-Pair-2001.nc /tmp/tp45e7e7cd_bd05_4714_a617_27c09cd269c2.nc /tmp/tpac79efaa_a6b2_4869_b047_62972be72429.nc\n",
			"Mon Sep 10 13:32:08 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2001.nc /tmp/tpf43628e7_83d0_4a16_bd5a_42915d7abb03.nc\n",
			"Thu Sep  6 10:40:07 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2001.nc\n",
			"Thu Sep  6 10:38:53 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2001_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2001.nc\n",
			"04-Oct-2017 17:51:47: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
