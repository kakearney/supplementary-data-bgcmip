netcdf CFS-atmos-northPacific-Tair-2018 {
dimensions:
	tair_time = UNLIMITED ; // (1451 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:missing_value = -1.e+34 ;
		Tair:_FillValue = -1.e+34 ;
		Tair:time = "tair_time" ;
		Tair:coordinates = "lon lat" ;
		Tair:height_above_ground = 2.f ;
		Tair:long_name = "surface air temperature" ;
		Tair:history = "From roms-cfs-atmos-Tair-2018" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double tair_time(tair_time) ;
		tair_time:units = "day since 1900-01-01 00:00:00" ;
		tair_time:time_origin = "01-JAN-1900 00:00:00" ;
		tair_time:axis = "T" ;
		tair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:23:27 2022: ncks -F -O -d tair_time,2,1452 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Tair-2018.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Tair-2018.nc\n",
			"Thu May 30 20:49:00 2019: Time overhang added\n",
			"Thu May 30 20:48:53 2019: ncrcat /tmp/tp04fcb445_371a_410b_b3ef_a56fc54dfaab.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Tair-2018.nc /tmp/tpb6993df0_74f5_43b7_a49e_f71b390ec57f.nc /tmp/tpf9a19502_b0bb_4e09_bedb_fa7c9710cfdd.nc\n",
			"Thu May 30 20:48:52 2019: ncks -F -d tair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Tair-2018.nc /tmp/tp04fcb445_371a_410b_b3ef_a56fc54dfaab.nc\n",
			"FERRET V7.4  29-May-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
