netcdf CFS-atmos-northPacific-Tair-1984 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:missing_value = -1.e+34 ;
		Tair:_FillValue = -1.e+34 ;
		Tair:time = "tair_time" ;
		Tair:coordinates = "lon lat" ;
		Tair:height_above_ground = 2.f ;
		Tair:long_name = "surface air temperature" ;
		Tair:history = "From roms-cfs-atmos-Tair-1984" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double tair_time(tair_time) ;
		tair_time:units = "day since 1900-01-01 00:00:00" ;
		tair_time:time_origin = "01-JAN-1900 00:00:00" ;
		tair_time:axis = "T" ;
		tair_time:standard_name = "time" ;

// global attributes:
		:history = "Thu Nov  3 15:34:31 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Tair-1984.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1984/CFS-atmos-northPacific-Tair-1984.nc\n",
			"Wed Nov 20 13:44:21 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:44:17 2019: ncrcat /tmp/tpbad993b8_cb06_4007_a57e_d934eb887db0.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Tair-1984.nc /tmp/tp99f1fad5_116c_4bd5_b936_fa913d57dc8c.nc /tmp/tpc40ce1a1_3952_4ffa_a5f3_f48e197b40a4.nc\n",
			"Wed Nov 20 13:44:14 2019: ncks -F -d tair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Tair-1984.nc /tmp/tpbad993b8_cb06_4007_a57e_d934eb887db0.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
