netcdf CFS-atmos-northPacific-rain-2007 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:54:48 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2007/roms-cfs-atmos-rain-2007.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2007/CFS-atmos-northPacific-rain-2007.nc\n",
			"Mon Sep 10 13:50:59 2018: Time overhang added\n",
			"Mon Sep 10 13:50:55 2018: ncrcat /tmp/tpe694e913_94b4_4583_b844_295bfce13dd1.nc frc/roms-cfs-atmos-rain-2007.nc /tmp/tp3269a233_cac8_4840_90ee_b330e976b8a2.nc /tmp/tp5f108db8_b679_41af_958b_1c5ca4a2cf03.nc\n",
			"Mon Sep 10 13:50:55 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2007.nc /tmp/tpe694e913_94b4_4583_b844_295bfce13dd1.nc\n",
			"Thu Sep  6 11:46:20 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2007_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2007.nc\n",
			"04-Oct-2017 18:07:08: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
