netcdf CFS-ocean-Bering10K-N30-bryocn-1990 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	xi_rho = 182 ;
	xi_u = 181 ;
	xi_v = 182 ;
	s_rho = 30 ;
	eta_rho = 258 ;
	eta_u = 258 ;
	eta_v = 257 ;
variables:
	double bry_time(bry_time) ;
		bry_time:standard_name = "time" ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:axis = "T" ;
	double zeta_south(bry_time, xi_rho) ;
		zeta_south:long_name = "free-surface, southern boundary condition" ;
		zeta_south:_FillValue = -999999. ;
		zeta_south:missing_value = -999999. ;
		zeta_south:unit = "meter" ;
		zeta_south:time = "bry_time" ;
		zeta_south:cell_methods = "bry_time: mean" ;
	double ubar_south(bry_time, xi_u) ;
		ubar_south:long_name = "vertically integrated u-momentum component, southern boundary condition" ;
		ubar_south:_FillValue = -999999. ;
		ubar_south:missing_value = -999999. ;
		ubar_south:unit = "meter second-1" ;
		ubar_south:time = "bry_time" ;
		ubar_south:cell_methods = "bry_time: mean" ;
	double vbar_south(bry_time, xi_v) ;
		vbar_south:long_name = "vertically integrated v-momentum component, southern boundary condition" ;
		vbar_south:_FillValue = -999999. ;
		vbar_south:missing_value = -999999. ;
		vbar_south:unit = "meter second-1" ;
		vbar_south:time = "bry_time" ;
		vbar_south:cell_methods = "bry_time: mean" ;
	double u_south(bry_time, s_rho, xi_u) ;
		u_south:long_name = "u-momentum component, southern boundary condition" ;
		u_south:_FillValue = -999999. ;
		u_south:missing_value = -999999. ;
		u_south:unit = "meter second-1" ;
		u_south:time = "bry_time" ;
		u_south:cell_methods = "bry_time: mean" ;
	double v_south(bry_time, s_rho, xi_v) ;
		v_south:long_name = "v-momentum component, southern boundary condition" ;
		v_south:_FillValue = -999999. ;
		v_south:missing_value = -999999. ;
		v_south:unit = "meter second-1" ;
		v_south:time = "bry_time" ;
		v_south:cell_methods = "bry_time: mean" ;
	double temp_south(bry_time, s_rho, xi_rho) ;
		temp_south:long_name = "potential temperature, southern boundary condition" ;
		temp_south:_FillValue = -999999. ;
		temp_south:missing_value = -999999. ;
		temp_south:unit = "Celsius" ;
		temp_south:time = "bry_time" ;
		temp_south:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:_FillValue = -999999. ;
		salt_south:missing_value = -999999. ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double zeta_west(bry_time, eta_rho) ;
		zeta_west:long_name = "free-surface, western boundary condition" ;
		zeta_west:_FillValue = -999999. ;
		zeta_west:missing_value = -999999. ;
		zeta_west:unit = "meter" ;
		zeta_west:time = "bry_time" ;
		zeta_west:cell_methods = "bry_time: mean" ;
	double ubar_west(bry_time, eta_u) ;
		ubar_west:long_name = "vertically integrated u-momentum component, western boundary condition" ;
		ubar_west:_FillValue = -999999. ;
		ubar_west:missing_value = -999999. ;
		ubar_west:unit = "meter second-1" ;
		ubar_west:time = "bry_time" ;
		ubar_west:cell_methods = "bry_time: mean" ;
	double vbar_west(bry_time, eta_v) ;
		vbar_west:long_name = "vertically integrated v-momentum component, western boundary condition" ;
		vbar_west:_FillValue = -999999. ;
		vbar_west:missing_value = -999999. ;
		vbar_west:unit = "meter second-1" ;
		vbar_west:time = "bry_time" ;
		vbar_west:cell_methods = "bry_time: mean" ;
	double u_west(bry_time, s_rho, eta_u) ;
		u_west:long_name = "u-momentum component, western boundary condition" ;
		u_west:_FillValue = -999999. ;
		u_west:missing_value = -999999. ;
		u_west:unit = "meter second-1" ;
		u_west:time = "bry_time" ;
		u_west:cell_methods = "bry_time: mean" ;
	double v_west(bry_time, s_rho, eta_v) ;
		v_west:long_name = "v-momentum component, western boundary condition" ;
		v_west:_FillValue = -999999. ;
		v_west:missing_value = -999999. ;
		v_west:unit = "meter second-1" ;
		v_west:time = "bry_time" ;
		v_west:cell_methods = "bry_time: mean" ;
	double temp_west(bry_time, s_rho, eta_rho) ;
		temp_west:long_name = "potential temperature, western boundary condition" ;
		temp_west:_FillValue = -999999. ;
		temp_west:missing_value = -999999. ;
		temp_west:unit = "Celsius" ;
		temp_west:time = "bry_time" ;
		temp_west:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:_FillValue = -999999. ;
		salt_west:missing_value = -999999. ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double zeta_east(bry_time, eta_rho) ;
		zeta_east:long_name = "free-surface, eastern boundary condition" ;
		zeta_east:_FillValue = -999999. ;
		zeta_east:missing_value = -999999. ;
		zeta_east:unit = "meter" ;
		zeta_east:time = "bry_time" ;
		zeta_east:cell_methods = "bry_time: mean" ;
	double ubar_east(bry_time, eta_u) ;
		ubar_east:long_name = "vertically integrated u-momentum component, eastern boundary condition" ;
		ubar_east:_FillValue = -999999. ;
		ubar_east:missing_value = -999999. ;
		ubar_east:unit = "meter second-1" ;
		ubar_east:time = "bry_time" ;
		ubar_east:cell_methods = "bry_time: mean" ;
	double vbar_east(bry_time, eta_v) ;
		vbar_east:long_name = "vertically integrated v-momentum component, eastern boundary condition" ;
		vbar_east:_FillValue = -999999. ;
		vbar_east:missing_value = -999999. ;
		vbar_east:unit = "meter second-1" ;
		vbar_east:time = "bry_time" ;
		vbar_east:cell_methods = "bry_time: mean" ;
	double u_east(bry_time, s_rho, eta_u) ;
		u_east:long_name = "u-momentum component, eastern boundary condition" ;
		u_east:_FillValue = -999999. ;
		u_east:missing_value = -999999. ;
		u_east:unit = "meter second-1" ;
		u_east:time = "bry_time" ;
		u_east:cell_methods = "bry_time: mean" ;
	double v_east(bry_time, s_rho, eta_v) ;
		v_east:long_name = "v-momentum component, eastern boundary condition" ;
		v_east:_FillValue = -999999. ;
		v_east:missing_value = -999999. ;
		v_east:unit = "meter second-1" ;
		v_east:time = "bry_time" ;
		v_east:cell_methods = "bry_time: mean" ;
	double temp_east(bry_time, s_rho, eta_rho) ;
		temp_east:long_name = "potential temperature, eastern boundary condition" ;
		temp_east:_FillValue = -999999. ;
		temp_east:missing_value = -999999. ;
		temp_east:unit = "Celsius" ;
		temp_east:time = "bry_time" ;
		temp_east:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:_FillValue = -999999. ;
		salt_east:missing_value = -999999. ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.1.0 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:type = "BOUNDARY file" ;
		:history = "Fri Sep 22 16:55:21 2023: cdo setmissval,-999999 CFS/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc test.nc\n",
			"Fri Sep 22 16:37:57 2023: cdo setmissval,nan CFS/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc test.nc\n",
			"Mon Dec 12 10:29:38 2022: ncrcat -O <>/final/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad73.nc <>/final/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc\n",
			"Fri Dec  9 16:24:34 2022: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad01.nc <>/final/1990/CFS-ocean-Bering10K-N30-bryocn-1990.nc\n",
			"Fri Dec  9 16:24:34 2022: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad01.nc\n",
			"Fri Dec  9 16:24:34 2022: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1990010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1990pentad01.nc\n",
			"Fri Dec 09 16:09:28 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
		:CDO = "Climate Data Operators version 2.1.0 (https://mpimet.mpg.de/cdo)" ;
}
