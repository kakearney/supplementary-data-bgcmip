netcdf CFS-atmos-northPacific-Pair-2010 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:00:01 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2010/roms-cfs-atmos-Pair-2010.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Pair-2010.nc\n",
			"Mon Sep 10 13:32:59 2018: Time overhang added\n",
			"Mon Sep 10 13:32:56 2018: ncrcat /tmp/tpd024e835_ad8d_45f4_8a0e_4d1bf6692df0.nc frc/roms-cfs-atmos-Pair-2010.nc /tmp/tp46110caf_242a_4269_b2b3_a56c6ca18719.nc /tmp/tp1775ca5c_940b_4e02_8428_2f8520ad0288.nc\n",
			"Mon Sep 10 13:32:56 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2010.nc /tmp/tpd024e835_ad8d_45f4_8a0e_4d1bf6692df0.nc\n",
			"Thu Sep  6 12:05:51 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2010.nc\n",
			"Thu Sep  6 12:04:59 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2010_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2010.nc\n",
			"04-Oct-2017 18:11:27: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
