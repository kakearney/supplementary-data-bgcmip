netcdf CFS-atmos-northPacific-swrad-2015 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:54:00 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2015/roms-cfs-atmos-swrad-2015.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-swrad-2015.nc\n",
			"Mon Sep 10 14:04:34 2018: Time overhang added\n",
			"Mon Sep 10 14:04:31 2018: ncrcat /tmp/tp3bc90838_d884_4d70_9570_dc05ebdba6ad.nc frc/roms-cfs-atmos-swrad-2015.nc /tmp/tp03185ee1_d718_401e_aeef_3e4c092df716.nc /tmp/tp7e5cc502_a1cd_4e54_8505_aa3119edfcd8.nc\n",
			"Mon Sep 10 14:04:31 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-2015.nc /tmp/tp3bc90838_d884_4d70_9570_dc05ebdba6ad.nc\n",
			"Thu Sep  6 13:52:39 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2015_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-2015.nc\n",
			"04-Oct-2017 18:30:57: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
