netcdf CFS-atmos-northPacific-Pair-2012 {
dimensions:
	pair_time = UNLIMITED ; // (1464 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:13:33 2022: ncks -F -O -d pair_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2012/roms-cfs-atmos-Pair-2012.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Pair-2012.nc\n",
			"Mon Sep 10 13:33:20 2018: Time overhang added\n",
			"Mon Sep 10 13:33:12 2018: ncrcat /tmp/tp396a0a60_c70b_4ec9_bc8b_70712599cf85.nc frc/roms-cfs-atmos-Pair-2012.nc /tmp/tp263637f7_2127_4b67_9786_d5b9c22facea.nc /tmp/tp8fd0b8f4_84e6_4043_be22_1171b03e755f.nc\n",
			"Mon Sep 10 13:33:12 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2012.nc /tmp/tp396a0a60_c70b_4ec9_bc8b_70712599cf85.nc\n",
			"Thu Sep  6 12:33:19 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2012.nc\n",
			"Thu Sep  6 12:31:44 2018: ncks -O -F -d air_time,2,1465 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2012_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2012.nc\n",
			"04-Oct-2017 18:17:20: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
