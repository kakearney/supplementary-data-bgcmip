netcdf CFS-atmos-northPacific-Uwind-1995 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:37:17 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1995/roms-cfs-atmos-Uwind-1995.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1995/CFS-atmos-northPacific-Uwind-1995.nc\n",
			"Mon Sep 10 13:40:23 2018: Time overhang added\n",
			"Mon Sep 10 13:40:20 2018: ncrcat /tmp/tp5a7ee844_f01b_41ba_ac27_12781fd1c6e3.nc frc/roms-cfs-atmos-Uwind-1995.nc /tmp/tpad934df3_5193_4ea9_bd41_3b767e070f77.nc /tmp/tp30cc00bd_99a7_4da3_94eb_b580f9b0f79c.nc\n",
			"Mon Sep 10 13:40:20 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-1995.nc /tmp/tp5a7ee844_f01b_41ba_ac27_12781fd1c6e3.nc\n",
			"Thu Sep  6 09:54:18 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1995_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-1995.nc\n",
			"04-Oct-2017 17:38:16: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
