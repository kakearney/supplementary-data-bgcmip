netcdf CFS-atmos-northPacific-swrad-1998 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:46:47 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1998/roms-cfs-atmos-swrad-1998.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1998/CFS-atmos-northPacific-swrad-1998.nc\n",
			"Mon Sep 10 14:03:47 2018: Time overhang added\n",
			"Mon Sep 10 14:03:45 2018: ncrcat /tmp/tpee5051cc_9e5f_4e36_86d9_9146108dc796.nc frc/roms-cfs-atmos-swrad-1998.nc /tmp/tpf7323256_4aa4_4d2e_9b1c_0c025eb834df.nc /tmp/tp1f2402ac_9c20_4e3c_9ff7_2bb034937457.nc\n",
			"Mon Sep 10 14:03:45 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-1998.nc /tmp/tpee5051cc_9e5f_4e36_86d9_9146108dc796.nc\n",
			"Thu Sep  6 10:18:06 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1998_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-1998.nc\n",
			"04-Oct-2017 17:45:31: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
