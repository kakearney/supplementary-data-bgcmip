netcdf CFS-atmos-northPacific-Pair-2002 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:03 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2002/roms-cfs-atmos-Pair-2002.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2002/CFS-atmos-northPacific-Pair-2002.nc\n",
			"Mon Sep 10 13:32:18 2018: Time overhang added\n",
			"Mon Sep 10 13:32:14 2018: ncrcat /tmp/tpf715df0b_0af9_4df7_b459_8fea8daf2bc2.nc frc/roms-cfs-atmos-Pair-2002.nc /tmp/tpb1f00d3b_26c0_48d6_a010_24da3aaa306e.nc /tmp/tp4141df56_5072_429b_86c6_0097bb5c4975.nc\n",
			"Mon Sep 10 13:32:14 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2002.nc /tmp/tpf715df0b_0af9_4df7_b459_8fea8daf2bc2.nc\n",
			"Thu Sep  6 10:50:15 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2002.nc\n",
			"Thu Sep  6 10:48:57 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2002_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2002.nc\n",
			"04-Oct-2017 17:54:31: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
