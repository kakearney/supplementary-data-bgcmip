netcdf CFS-atmos-northPacific-lwrad-2010 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:02:04 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2010/roms-cfs-atmos-lwrad-2010.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-lwrad-2010.nc\n",
			"Mon Sep 10 13:47:56 2018: Time overhang added\n",
			"Mon Sep 10 13:47:52 2018: ncrcat /tmp/tp7fa00668_bb2e_4812_8ed7_0efb193e8820.nc frc/roms-cfs-atmos-lwrad-2010.nc /tmp/tpbfef04a8_abeb_4bd3_8594_6a21b0f62015.nc /tmp/tpbe1a10cb_f054_4dae_9064_cda49d41c280.nc\n",
			"Mon Sep 10 13:47:52 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2010.nc /tmp/tp7fa00668_bb2e_4812_8ed7_0efb193e8820.nc\n",
			"Thu Sep  6 12:09:23 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2010_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2010.nc\n",
			"04-Oct-2017 18:12:10: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
