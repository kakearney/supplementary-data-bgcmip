netcdf CFS-atmos-northPacific-Tair-2002 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:16 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2002/roms-cfs-atmos-Tair-2002.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2002/CFS-atmos-northPacific-Tair-2002.nc\n",
			"Mon Sep 10 13:38:07 2018: Time overhang added\n",
			"Mon Sep 10 13:38:03 2018: ncrcat /tmp/tp7e7b2da1_5e68_4203_ac06_4bc829ffc735.nc frc/roms-cfs-atmos-Tair-2002.nc /tmp/tpb6b18593_e461_4139_8322_7c78d73a8889.nc /tmp/tp55166155_3a3f_4d6f_901f_de1f32045811.nc\n",
			"Mon Sep 10 13:38:03 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2002.nc /tmp/tp7e7b2da1_5e68_4203_ac06_4bc829ffc735.nc\n",
			"Thu Sep  6 10:52:06 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2002.nc\n",
			"Thu Sep  6 10:50:57 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2002_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2002.nc\n",
			"04-Oct-2017 17:54:31: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
