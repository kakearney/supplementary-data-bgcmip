netcdf CFS-atmos-northPacific-rain-2010 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:02:10 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2010/roms-cfs-atmos-rain-2010.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-rain-2010.nc\n",
			"Mon Sep 10 13:51:16 2018: Time overhang added\n",
			"Mon Sep 10 13:51:12 2018: ncrcat /tmp/tp1378c121_b24d_4207_a540_f1210b34b879.nc frc/roms-cfs-atmos-rain-2010.nc /tmp/tp624e437e_3564_403c_9b4c_a6ff0f3ac8a5.nc /tmp/tp916e0c34_c41b_4f04_b597_6894c316bc89.nc\n",
			"Mon Sep 10 13:51:12 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2010.nc /tmp/tp1378c121_b24d_4207_a540_f1210b34b879.nc\n",
			"Thu Sep  6 12:10:03 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2010_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2010.nc\n",
			"04-Oct-2017 18:13:08: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
