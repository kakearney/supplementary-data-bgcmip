netcdf CFS-atmos-northPacific-rain-2016 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	rain_time = UNLIMITED ; // (1448 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Mon Oct 31 12:06:21 2022: ncks -F -O -d rain_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2016/roms-cfs-atmos-rain-2016.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-rain-2016.nc\n",
			"Mon Sep 10 14:03:14 2018: Time overhang added\n",
			"Mon Sep 10 14:03:06 2018: ncrcat /tmp/tp01eea2e5_b7b5_4c9c_b410_59c11b25a51e.nc frc/roms-cfs-atmos-rain-2016.nc /tmp/tpc470876b_8566_41ad_a762_cb9fb3a24a2e.nc /tmp/tpcdb7a19f_730c_4af1_999f_2daa2ad87860.nc\n",
			"Mon Sep 10 14:03:06 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2016.nc /tmp/tp01eea2e5_b7b5_4c9c_b410_59c11b25a51e.nc\n",
			"Thu Sep  6 14:15:29 2018: ncks -O -F -d rain_time,2,1449 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2016_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2016.nc\n",
			"04-Oct-2017 18:35:56: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
