netcdf CFS-atmos-northPacific-Pair-1994 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:missing_value = -1.e+34 ;
		Pair:_FillValue = -1.e+34 ;
		Pair:time = "pair_time" ;
		Pair:coordinates = "lon lat" ;
		Pair:long_name = "atmos pressure" ;
		Pair:history = "From roms-cfs-atmos-Pair-1994" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double pair_time(pair_time) ;
		pair_time:units = "day since 1900-01-01 00:00:00" ;
		pair_time:time_origin = "01-JAN-1900 00:00:00" ;
		pair_time:axis = "T" ;
		pair_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:34:20 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1994/roms-cfs-atmos-Pair-1994.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1994/CFS-atmos-northPacific-Pair-1994.nc\n",
			"Wed Nov 20 14:04:39 2019: Time overhang added to both ends\n",
			"Wed Nov 20 14:04:33 2019: ncrcat /tmp/tp46291be2_c8a3_424c_b755_9236086a642b.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1994/roms-cfs-atmos-Pair-1994.nc /tmp/tp2f8cb788_4aad_46ff_8234_cfbb2e5f8d7e.nc /tmp/tpfb07ae02_04b6_4d91_80b8_b38265b2c790.nc\n",
			"Wed Nov 20 14:04:31 2019: ncks -F -d pair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1994/roms-cfs-atmos-Pair-1994.nc /tmp/tp46291be2_c8a3_424c_b755_9236086a642b.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
