netcdf CFS-atmos-northPacific-Vwind-2001 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:50:00 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2001/roms-cfs-atmos-Vwind-2001.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2001/CFS-atmos-northPacific-Vwind-2001.nc\n",
			"Mon Sep 10 13:44:01 2018: Time overhang added\n",
			"Mon Sep 10 13:43:57 2018: ncrcat /tmp/tp90834b25_072b_4aed_bc89_2f6ca22aff2b.nc frc/roms-cfs-atmos-Vwind-2001.nc /tmp/tp846065a5_2106_43f4_82a0_17285ea89edb.nc /tmp/tp7c41c271_be8c_438f_a9ed_ca4c815d2b56.nc\n",
			"Mon Sep 10 13:43:57 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2001.nc /tmp/tp90834b25_072b_4aed_bc89_2f6ca22aff2b.nc\n",
			"Thu Sep  6 10:47:48 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2001_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2001.nc\n",
			"04-Oct-2017 17:53:12: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
