netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-1997 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:01:33 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 14:58:43 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1997/CFS-ocean-NEP-N30-bryocn-1997.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1997/CFS-ocean-ESPER-NEP-N30-brycarbon-1997.nc\n",
			"Sat Dec 17 02:34:23 2022: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad73.nc <>/final/1997/CFS-ocean-NEP-N30-bryocn-1997.nc\n",
			"Sat Dec 17 02:33:02 2022: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad01.nc\n",
			"Sat Dec 17 02:33:01 2022: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1997010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1997pentad01.nc\n",
			"Fri Dec 16 19:03:06 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
