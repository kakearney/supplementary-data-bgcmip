netcdf CFS-atmos-northPacific-Vwind-2019 {
dimensions:
	wind_time = UNLIMITED ; // (1457 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:missing_value = -1.e+34 ;
		Vwind:_FillValue = -1.e+34 ;
		Vwind:time = "wind_time" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:height_above_ground1 = 10.f ;
		Vwind:long_name = "V wind" ;
		Vwind:history = "From roms-cfs-atmos-Vwind-2019" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:39:35 2022: ncks -F -O -d wind_time,2,1458 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Vwind-2019.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Vwind-2019.nc\n",
			"Fri Mar 27 16:04:34 2020: Time overhang added to both ends\n",
			"Fri Mar 27 16:04:25 2020: ncrcat /tmp/tp915cee76_4277_4113_894d_439887c43e3c.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Vwind-2019.nc /tmp/tp0b941097_ed94_4331_a1d8_9096fcec43dd.nc /tmp/tp4cd1322c_6ef4_45a9_b117_65d6ffbf93ba.nc\n",
			"Fri Mar 27 16:04:23 2020: ncks -F -d wind_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Vwind-2019.nc /tmp/tp915cee76_4277_4113_894d_439887c43e3c.nc\n",
			"FERRET V7.4   4-Mar-20" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
