netcdf CFS-ocean-NEP-N30-bryocn-2020 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	eta_rho = 642 ;
	s_rho = 30 ;
	xi_rho = 226 ;
	eta_u = 642 ;
	xi_u = 225 ;
	eta_v = 641 ;
	xi_v = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:standard_name = "time" ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:axis = "T" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:_FillValue = -999999. ;
		salt_east:missing_value = -999999. ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:_FillValue = -999999. ;
		salt_south:missing_value = -999999. ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:_FillValue = -999999. ;
		salt_west:missing_value = -999999. ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double temp_east(bry_time, s_rho, eta_rho) ;
		temp_east:long_name = "potential temperature, eastern boundary condition" ;
		temp_east:_FillValue = -999999. ;
		temp_east:missing_value = -999999. ;
		temp_east:unit = "Celsius" ;
		temp_east:time = "bry_time" ;
		temp_east:cell_methods = "bry_time: mean" ;
	double temp_south(bry_time, s_rho, xi_rho) ;
		temp_south:long_name = "potential temperature, southern boundary condition" ;
		temp_south:_FillValue = -999999. ;
		temp_south:missing_value = -999999. ;
		temp_south:unit = "Celsius" ;
		temp_south:time = "bry_time" ;
		temp_south:cell_methods = "bry_time: mean" ;
	double temp_west(bry_time, s_rho, eta_rho) ;
		temp_west:long_name = "potential temperature, western boundary condition" ;
		temp_west:_FillValue = -999999. ;
		temp_west:missing_value = -999999. ;
		temp_west:unit = "Celsius" ;
		temp_west:time = "bry_time" ;
		temp_west:cell_methods = "bry_time: mean" ;
	double u_east(bry_time, s_rho, eta_u) ;
		u_east:long_name = "u-momentum component, eastern boundary condition" ;
		u_east:_FillValue = -999999. ;
		u_east:missing_value = -999999. ;
		u_east:unit = "meter second-1" ;
		u_east:time = "bry_time" ;
		u_east:cell_methods = "bry_time: mean" ;
	double u_south(bry_time, s_rho, xi_u) ;
		u_south:long_name = "u-momentum component, southern boundary condition" ;
		u_south:_FillValue = -999999. ;
		u_south:missing_value = -999999. ;
		u_south:unit = "meter second-1" ;
		u_south:time = "bry_time" ;
		u_south:cell_methods = "bry_time: mean" ;
	double u_west(bry_time, s_rho, eta_u) ;
		u_west:long_name = "u-momentum component, western boundary condition" ;
		u_west:_FillValue = -999999. ;
		u_west:missing_value = -999999. ;
		u_west:unit = "meter second-1" ;
		u_west:time = "bry_time" ;
		u_west:cell_methods = "bry_time: mean" ;
	double ubar_east(bry_time, eta_u) ;
		ubar_east:long_name = "vertically integrated u-momentum component, eastern boundary condition" ;
		ubar_east:_FillValue = -999999. ;
		ubar_east:missing_value = -999999. ;
		ubar_east:unit = "meter second-1" ;
		ubar_east:time = "bry_time" ;
		ubar_east:cell_methods = "bry_time: mean" ;
	double ubar_south(bry_time, xi_u) ;
		ubar_south:long_name = "vertically integrated u-momentum component, southern boundary condition" ;
		ubar_south:_FillValue = -999999. ;
		ubar_south:missing_value = -999999. ;
		ubar_south:unit = "meter second-1" ;
		ubar_south:time = "bry_time" ;
		ubar_south:cell_methods = "bry_time: mean" ;
	double ubar_west(bry_time, eta_u) ;
		ubar_west:long_name = "vertically integrated u-momentum component, western boundary condition" ;
		ubar_west:_FillValue = -999999. ;
		ubar_west:missing_value = -999999. ;
		ubar_west:unit = "meter second-1" ;
		ubar_west:time = "bry_time" ;
		ubar_west:cell_methods = "bry_time: mean" ;
	double v_east(bry_time, s_rho, eta_v) ;
		v_east:long_name = "v-momentum component, eastern boundary condition" ;
		v_east:_FillValue = -999999. ;
		v_east:missing_value = -999999. ;
		v_east:unit = "meter second-1" ;
		v_east:time = "bry_time" ;
		v_east:cell_methods = "bry_time: mean" ;
	double v_south(bry_time, s_rho, xi_v) ;
		v_south:long_name = "v-momentum component, southern boundary condition" ;
		v_south:_FillValue = -999999. ;
		v_south:missing_value = -999999. ;
		v_south:unit = "meter second-1" ;
		v_south:time = "bry_time" ;
		v_south:cell_methods = "bry_time: mean" ;
	double v_west(bry_time, s_rho, eta_v) ;
		v_west:long_name = "v-momentum component, western boundary condition" ;
		v_west:_FillValue = -999999. ;
		v_west:missing_value = -999999. ;
		v_west:unit = "meter second-1" ;
		v_west:time = "bry_time" ;
		v_west:cell_methods = "bry_time: mean" ;
	double vbar_east(bry_time, eta_v) ;
		vbar_east:long_name = "vertically integrated v-momentum component, eastern boundary condition" ;
		vbar_east:_FillValue = -999999. ;
		vbar_east:missing_value = -999999. ;
		vbar_east:unit = "meter second-1" ;
		vbar_east:time = "bry_time" ;
		vbar_east:cell_methods = "bry_time: mean" ;
	double vbar_south(bry_time, xi_v) ;
		vbar_south:long_name = "vertically integrated v-momentum component, southern boundary condition" ;
		vbar_south:_FillValue = -999999. ;
		vbar_south:missing_value = -999999. ;
		vbar_south:unit = "meter second-1" ;
		vbar_south:time = "bry_time" ;
		vbar_south:cell_methods = "bry_time: mean" ;
	double vbar_west(bry_time, eta_v) ;
		vbar_west:long_name = "vertically integrated v-momentum component, western boundary condition" ;
		vbar_west:_FillValue = -999999. ;
		vbar_west:missing_value = -999999. ;
		vbar_west:unit = "meter second-1" ;
		vbar_west:time = "bry_time" ;
		vbar_west:cell_methods = "bry_time: mean" ;
	double zeta_east(bry_time, eta_rho) ;
		zeta_east:long_name = "free-surface, eastern boundary condition" ;
		zeta_east:_FillValue = -999999. ;
		zeta_east:missing_value = -999999. ;
		zeta_east:unit = "meter" ;
		zeta_east:time = "bry_time" ;
		zeta_east:cell_methods = "bry_time: mean" ;
	double zeta_south(bry_time, xi_rho) ;
		zeta_south:long_name = "free-surface, southern boundary condition" ;
		zeta_south:_FillValue = -999999. ;
		zeta_south:missing_value = -999999. ;
		zeta_south:unit = "meter" ;
		zeta_south:time = "bry_time" ;
		zeta_south:cell_methods = "bry_time: mean" ;
	double zeta_west(bry_time, eta_rho) ;
		zeta_west:long_name = "free-surface, western boundary condition" ;
		zeta_west:_FillValue = -999999. ;
		zeta_west:missing_value = -999999. ;
		zeta_west:unit = "meter" ;
		zeta_west:time = "bry_time" ;
		zeta_west:cell_methods = "bry_time: mean" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.1.0 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:type = "BOUNDARY file" ;
		:history = "Fri Sep 22 16:55:49 2023: cdo setmissval,-999999 CFS/2020/CFS-ocean-NEP-N30-bryocn-2020.nc test.nc\n",
			"Fri Sep 22 16:38:37 2023: cdo setmissval,nan CFS/2020/CFS-ocean-NEP-N30-bryocn-2020.nc test.nc\n",
			"Thu Jan 12 22:09:32 2023: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad73.nc <>/final/2020/CFS-ocean-NEP-N30-bryocn-2020.nc\n",
			"Thu Jan 12 22:02:58 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad01.nc\n",
			"Thu Jan 12 22:02:57 2023: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad01.nc\n",
			"Thu Jan 12 22:02:55 2023: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2020010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2020pentad01.nc\n",
			"Thu Jan 12 08:15:15 2023: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
		:CDO = "Climate Data Operators version 2.1.0 (https://mpimet.mpg.de/cdo)" ;
}
