netcdf INIbgc_BEST_NPZ_NEP {
dimensions:
	xi_rho = 226 ;
	eta_rho = 642 ;
	s_rho = 30 ;
	benlayer = 1 ;
	ocean_time = UNLIMITED ; // (1 currently)
variables:
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 1900-01-01 00:00:00" ;
		ocean_time:calendar = "standard" ;
	double NO3(ocean_time, s_rho, eta_rho, xi_rho) ;
		NO3:long_name = "Nitrate concentration" ;
		NO3:unit = "mmol N m^-3" ;
		NO3:time = "ocean_time" ;
		NO3:_FillValue = 1.e+36 ;
	double NH4(ocean_time, s_rho, eta_rho, xi_rho) ;
		NH4:long_name = "Ammonium concentration" ;
		NH4:unit = "mmol N m^-3" ;
		NH4:time = "ocean_time" ;
		NH4:_FillValue = 1.e+36 ;
	double PhS(ocean_time, s_rho, eta_rho, xi_rho) ;
		PhS:long_name = "Small phytoplankton concentration" ;
		PhS:unit = "mg C m^-3" ;
		PhS:time = "ocean_time" ;
		PhS:_FillValue = 1.e+36 ;
	double PhL(ocean_time, s_rho, eta_rho, xi_rho) ;
		PhL:long_name = "Large phytoplankton concentration" ;
		PhL:unit = "mg C m^-3" ;
		PhL:time = "ocean_time" ;
		PhL:_FillValue = 1.e+36 ;
	double MZL(ocean_time, s_rho, eta_rho, xi_rho) ;
		MZL:long_name = "Microzooplankton concentration" ;
		MZL:unit = "mg C m^-3" ;
		MZL:time = "ocean_time" ;
		MZL:_FillValue = 1.e+36 ;
	double Cop(ocean_time, s_rho, eta_rho, xi_rho) ;
		Cop:long_name = "Small copepod concentration" ;
		Cop:unit = "mg C m^-3" ;
		Cop:time = "ocean_time" ;
		Cop:_FillValue = 1.e+36 ;
	double NCaS(ocean_time, s_rho, eta_rho, xi_rho) ;
		NCaS:long_name = "On-shelf large copepod concentration" ;
		NCaS:unit = "mg C m^-3" ;
		NCaS:time = "ocean_time" ;
		NCaS:_FillValue = 1.e+36 ;
	double EupS(ocean_time, s_rho, eta_rho, xi_rho) ;
		EupS:long_name = "On-shelf euphausiid concentration" ;
		EupS:unit = "mg C m^-3" ;
		EupS:time = "ocean_time" ;
		EupS:_FillValue = 1.e+36 ;
	double NCaO(ocean_time, s_rho, eta_rho, xi_rho) ;
		NCaO:long_name = "Offshore large copepod concentration" ;
		NCaO:unit = "mg C m^-3" ;
		NCaO:time = "ocean_time" ;
		NCaO:_FillValue = 1.e+36 ;
	double EupO(ocean_time, s_rho, eta_rho, xi_rho) ;
		EupO:long_name = "Offshore euphausiid concentration" ;
		EupO:unit = "mg C m^-3" ;
		EupO:time = "ocean_time" ;
		EupO:_FillValue = 1.e+36 ;
	double Det(ocean_time, s_rho, eta_rho, xi_rho) ;
		Det:long_name = "Slow-sinking detritus concentration" ;
		Det:unit = "mg C m^-3" ;
		Det:time = "ocean_time" ;
		Det:_FillValue = 1.e+36 ;
	double DetF(ocean_time, s_rho, eta_rho, xi_rho) ;
		DetF:long_name = "Fast-sinking detritus concentration" ;
		DetF:unit = "mg C m^-3" ;
		DetF:time = "ocean_time" ;
		DetF:_FillValue = 1.e+36 ;
	double Jel(ocean_time, s_rho, eta_rho, xi_rho) ;
		Jel:long_name = "Jellyfish concentration" ;
		Jel:unit = "mg C m^-3" ;
		Jel:time = "ocean_time" ;
		Jel:_FillValue = 1.e+36 ;
	double Ben(ocean_time, benlayer, eta_rho, xi_rho) ;
		Ben:long_name = "Benthic infauna concentration" ;
		Ben:unit = "mg C m^-2" ;
		Ben:time = "ocean_time" ;
		Ben:_FillValue = 1.e+36 ;
	double DetBen(ocean_time, benlayer, eta_rho, xi_rho) ;
		DetBen:long_name = "Benthic detritus concentration" ;
		DetBen:unit = "mg C m^-2" ;
		DetBen:time = "ocean_time" ;
		DetBen:_FillValue = 1.e+36 ;
	double IcePhL(ocean_time, eta_rho, xi_rho) ;
		IcePhL:long_name = "Ice algae concentration" ;
		IcePhL:unit = "mg C m^-3" ;
		IcePhL:time = "ocean_time" ;
		IcePhL:_FillValue = 1.e+36 ;
	double IceNO3(ocean_time, eta_rho, xi_rho) ;
		IceNO3:long_name = "Ice nitrate concentration" ;
		IceNO3:unit = "mmol N m^-3" ;
		IceNO3:time = "ocean_time" ;
		IceNO3:_FillValue = 1.e+36 ;
	double IceNH4(ocean_time, eta_rho, xi_rho) ;
		IceNH4:long_name = "Ice ammonium concentration" ;
		IceNH4:unit = "mmol N m^-3" ;
		IceNH4:time = "ocean_time" ;
		IceNH4:_FillValue = 1.e+36 ;
	double Fe(ocean_time, s_rho, eta_rho, xi_rho) ;
		Fe:long_name = "Iron concentration" ;
		Fe:unit = "umol Fe m^-3" ;
		Fe:time = "ocean_time" ;
		Fe:_FillValue = 1.e+36 ;
	double alkalinity(ocean_time, s_rho, eta_rho, xi_rho) ;
		alkalinity:long_name = "total alkalinity" ;
		alkalinity:unit = "mmol C m^-3" ;
		alkalinity:time = "ocean_time" ;
		alkalinity:_FillValue = 1.e+36 ;
	double TIC(ocean_time, s_rho, eta_rho, xi_rho) ;
		TIC:long_name = "total inorganic carbon" ;
		TIC:unit = "mmol C m^-3" ;
		TIC:time = "ocean_time" ;
		TIC:_FillValue = 1.e+36 ;
	double oxygen(ocean_time, s_rho, eta_rho, xi_rho) ;
		oxygen:long_name = "dissolved oxygen concentration" ;
		oxygen:unit = "mmol O m^-3" ;
		oxygen:time = "ocean_time" ;
		oxygen:_FillValue = 1.e+36 ;

// global attributes:
		:type = "INITIALIZATION file" ;
		:history = "Wed Jan 25 11:27:09 2023: BGC data added: NO3, PO4, Alk, TIC, O2, SiO4: GLODAPv2.2016b Mapped Climatologies; Fe: Huang et al., 2022 climatology + GOANPZ analytical; Hfree, CO3: GLODAPv2 + CO2sys; producers/consumers: seed value; others: 0\n",
			"Wed Jan 25 11:27:07 2023: File schema created via ini_schema.m" ;
}
