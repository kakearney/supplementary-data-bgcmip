netcdf CFS-atmos-northPacific-lwrad-2003 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:17:22 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2003/roms-cfs-atmos-lwrad-2003.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2003/CFS-atmos-northPacific-lwrad-2003.nc\n",
			"Mon Sep 10 13:47:16 2018: Time overhang added\n",
			"Mon Sep 10 13:47:13 2018: ncrcat /tmp/tp94d450b3_19cd_4bb4_8107_fd9299919538.nc frc/roms-cfs-atmos-lwrad-2003.nc /tmp/tp3c0a31c4_4d10_4751_ab23_4ab5bba557dc.nc /tmp/tpe82edfc7_09a6_40cf_bfde_c5ca8f340586.nc\n",
			"Mon Sep 10 13:47:12 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2003.nc /tmp/tp94d450b3_19cd_4bb4_8107_fd9299919538.nc\n",
			"Thu Sep  6 11:03:54 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2003_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2003.nc\n",
			"04-Oct-2017 17:57:59: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
