netcdf CFS-atmos-northPacific-Vwind-1986 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:missing_value = -1.e+34 ;
		Vwind:_FillValue = -1.e+34 ;
		Vwind:time = "wind_time" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:height_above_ground1 = 10.f ;
		Vwind:long_name = "V wind" ;
		Vwind:history = "From roms-cfs-atmos-Vwind-1986" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:19:50 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-Vwind-1986.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1986/CFS-atmos-northPacific-Vwind-1986.nc\n",
			"Wed Nov 20 13:48:46 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:48:40 2019: ncrcat /tmp/tpde074e43_433b_4c5b_93f3_577efa69e4ac.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-Vwind-1986.nc /tmp/tp4bac0d19_03c9_4505_a1ff_056d66f288ac.nc /tmp/tpf1df6981_6cbe_41c0_b233_d9bf84d3f51d.nc\n",
			"Wed Nov 20 13:48:38 2019: ncks -F -d wind_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-Vwind-1986.nc /tmp/tpde074e43_433b_4c5b_93f3_577efa69e4ac.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
