netcdf CFS-atmos-northPacific-Qair-2008 {
dimensions:
	qair_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:55:53 2022: ncks -F -O -d qair_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2008/roms-cfs-atmos-Qair-2008.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2008/CFS-atmos-northPacific-Qair-2008.nc\n",
			"Mon Sep 10 13:35:44 2018: Time overhang added\n",
			"Mon Sep 10 13:35:40 2018: ncrcat /tmp/tp87df5560_cb8b_422d_b39b_4c19411f85eb.nc frc/roms-cfs-atmos-Qair-2008.nc /tmp/tp596cb4f1_3172_4f34_b6f0_f20893fdafd5.nc /tmp/tp3882423c_615c_499f_9270_8b2f060adb1d.nc\n",
			"Mon Sep 10 13:35:39 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2008.nc /tmp/tp87df5560_cb8b_422d_b39b_4c19411f85eb.nc\n",
			"Thu Sep  6 11:53:42 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2008.nc\n",
			"Thu Sep  6 11:53:00 2018: ncks -O -F -d air_time,2,1465 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2008_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2008.nc\n",
			"04-Oct-2017 18:07:27: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
