netcdf CFS-atmos-northPacific-swrad-2007 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:55:04 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2007/roms-cfs-atmos-swrad-2007.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2007/CFS-atmos-northPacific-swrad-2007.nc\n",
			"Mon Sep 10 14:04:06 2018: Time overhang added\n",
			"Mon Sep 10 14:04:05 2018: ncrcat /tmp/tp0330518b_784d_4e39_ab04_cd599e89e1c7.nc frc/roms-cfs-atmos-swrad-2007.nc /tmp/tp3337f653_3dc5_4367_8f1e_8e6320ac2b08.nc /tmp/tpcbc0b752_b31c_4c11_aabc_4bcc9e641658.nc\n",
			"Mon Sep 10 14:04:05 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-2007.nc /tmp/tp0330518b_784d_4e39_ab04_cd599e89e1c7.nc\n",
			"Thu Sep  6 11:47:08 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2007_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-2007.nc\n",
			"04-Oct-2017 18:06:26: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
