netcdf CFS-atmos-northPacific-Vwind-1996 {
dimensions:
	wind_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:42:25 2022: ncks -F -O -d wind_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1996/roms-cfs-atmos-Vwind-1996.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1996/CFS-atmos-northPacific-Vwind-1996.nc\n",
			"Mon Sep 10 13:43:33 2018: Time overhang added\n",
			"Mon Sep 10 13:43:29 2018: ncrcat /tmp/tp49de1d5f_46a1_4631_8f56_2ca53f706be3.nc frc/roms-cfs-atmos-Vwind-1996.nc /tmp/tp5d81f1ad_697b_4d1e_92f5_1bc9f645ee73.nc /tmp/tpb88e9509_aa4c_41d7_98c2_b93487668f49.nc\n",
			"Mon Sep 10 13:43:28 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-1996.nc /tmp/tp49de1d5f_46a1_4631_8f56_2ca53f706be3.nc\n",
			"Thu Sep  6 10:02:06 2018: ncks -O -F -d wind_time,2,1465 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1996_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-1996.nc\n",
			"04-Oct-2017 17:40:44: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
