netcdf CFS-atmos-northPacific-lwrad-2016 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	lrf_time = UNLIMITED ; // (1448 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Mon Oct 31 11:57:35 2022: ncks -F -O -d lrf_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2016/roms-cfs-atmos-lwrad-2016.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-lwrad-2016.nc\n",
			"Mon Sep 10 13:49:07 2018: Time overhang added\n",
			"Mon Sep 10 13:48:59 2018: ncrcat /tmp/tp71dbebc1_9f2f_473f_a873_77fe17b5a3fb.nc frc/roms-cfs-atmos-lwrad-2016.nc /tmp/tpfc14b7b8_30da_4722_a7f7_fe18cea27638.nc /tmp/tpc9b6091d_862f_4188_a7e6_e0acec9e40c2.nc\n",
			"Mon Sep 10 13:48:58 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2016.nc /tmp/tp71dbebc1_9f2f_473f_a873_77fe17b5a3fb.nc\n",
			"Thu Sep  6 14:14:18 2018: ncks -O -F -d lrf_time,2,1449 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2016_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2016.nc\n",
			"04-Oct-2017 18:34:12: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
