netcdf CFS-atmos-northPacific-rain-2009 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:59:52 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2009/roms-cfs-atmos-rain-2009.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-rain-2009.nc\n",
			"Mon Sep 10 13:51:10 2018: Time overhang added\n",
			"Mon Sep 10 13:51:06 2018: ncrcat /tmp/tp31b30f61_11d6_4d9f_bee0_15f656eca366.nc frc/roms-cfs-atmos-rain-2009.nc /tmp/tp29f35fbe_8783_4bc1_a013_68815187cc2c.nc /tmp/tp89da2408_543e_4b56_8c9c_a6e85a7c5f77.nc\n",
			"Mon Sep 10 13:51:06 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2009.nc /tmp/tp31b30f61_11d6_4d9f_bee0_15f656eca366.nc\n",
			"Thu Sep  6 12:02:35 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2009_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2009.nc\n",
			"04-Oct-2017 18:11:09: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
