netcdf CFS-atmos-northPacific-Vwind-1998 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:46:27 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1998/roms-cfs-atmos-Vwind-1998.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1998/CFS-atmos-northPacific-Vwind-1998.nc\n",
			"Mon Sep 10 13:43:44 2018: Time overhang added\n",
			"Mon Sep 10 13:43:41 2018: ncrcat /tmp/tpb2c356d8_88b7_4e2a_aaac_ce11cb45982d.nc frc/roms-cfs-atmos-Vwind-1998.nc /tmp/tp5d9df894_3313_4e12_bd49_3bf42acce67a.nc /tmp/tp08d8871b_7569_4164_8c81_422e362bdfe0.nc\n",
			"Mon Sep 10 13:43:40 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-1998.nc /tmp/tpb2c356d8_88b7_4e2a_aaac_ce11cb45982d.nc\n",
			"Thu Sep  6 10:19:15 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1998_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-1998.nc\n",
			"04-Oct-2017 17:45:35: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
