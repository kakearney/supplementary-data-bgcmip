netcdf ini_hindcastloop2_BEST_NPZ {
dimensions:
	ocean_time = UNLIMITED ; // (1 currently)
	s_w = 31 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
	tracer = 19 ;
	benlayer = 1 ;
	s_rho = 30 ;
	boundary = 4 ;
	eta_u = 258 ;
	xi_u = 181 ;
	eta_v = 257 ;
	xi_v = 182 ;
variables:
	float AKs(ocean_time, s_w, eta_rho, xi_rho) ;
		AKs:long_name = "salinity vertical diffusion coefficient" ;
		AKs:units = "meter2 second-1" ;
		AKs:time = "ocean_time" ;
		AKs:grid = "grid" ;
		AKs:location = "face" ;
		AKs:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKs:field = "AKs, scalar, series" ;
	float AKt(ocean_time, s_w, eta_rho, xi_rho) ;
		AKt:long_name = "temperature vertical diffusion coefficient" ;
		AKt:units = "meter2 second-1" ;
		AKt:time = "ocean_time" ;
		AKt:grid = "grid" ;
		AKt:location = "face" ;
		AKt:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKt:field = "AKt, scalar, series" ;
	float AKv(ocean_time, s_w, eta_rho, xi_rho) ;
		AKv:long_name = "vertical viscosity coefficient" ;
		AKv:units = "meter2 second-1" ;
		AKv:time = "ocean_time" ;
		AKv:grid = "grid" ;
		AKv:location = "face" ;
		AKv:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKv:field = "AKv, scalar, series" ;
	double Akt_bak(tracer) ;
		Akt_bak:long_name = "background vertical mixing coefficient for tracers" ;
		Akt_bak:units = "meter2 second-1" ;
	double Akv_bak ;
		Akv_bak:long_name = "background vertical mixing coefficient for momentum" ;
		Akv_bak:units = "meter2 second-1" ;
	float Ben(ocean_time, benlayer, eta_rho, xi_rho) ;
		Ben:long_name = "Benthic infauna concentration" ;
		Ben:units = "mg C m^-2" ;
		Ben:time = "ocean_time" ;
		Ben:grid = "grid" ;
		Ben:location = "face" ;
		Ben:coordinates = "lon_rho lat_rho benlayer ocean_time" ;
		Ben:field = "benthos, scalar, series" ;
		Ben:_FillValue = 1.e+37f ;
	double BenPred ;
		BenPred:long_name = "Quadratic mortality rate due to undefined predation" ;
		BenPred:units = "1/mgC/d" ;
	int BioIter ;
		BioIter:long_name = "number of iterations to achieve convergence" ;
	float Cop(ocean_time, s_rho, eta_rho, xi_rho) ;
		Cop:long_name = "Small copepod concentration" ;
		Cop:units = "mg C m^-3" ;
		Cop:time = "ocean_time" ;
		Cop:grid = "grid" ;
		Cop:location = "face" ;
		Cop:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		Cop:field = "copepod, scalar, series" ;
		Cop:_FillValue = 1.e+37f ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
		Cs_r:field = "Cs_r, scalar" ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
		Cs_w:field = "Cs_w, scalar" ;
	float Det(ocean_time, s_rho, eta_rho, xi_rho) ;
		Det:long_name = "Slow-sinking detritus concentration" ;
		Det:units = "mg C m^-3" ;
		Det:time = "ocean_time" ;
		Det:grid = "grid" ;
		Det:location = "face" ;
		Det:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		Det:field = "detritus, scalar, series" ;
		Det:_FillValue = 1.e+37f ;
	float DetBen(ocean_time, benlayer, eta_rho, xi_rho) ;
		DetBen:long_name = "Benthic detritus concentration" ;
		DetBen:units = "mg C m^-2" ;
		DetBen:time = "ocean_time" ;
		DetBen:grid = "grid" ;
		DetBen:location = "face" ;
		DetBen:coordinates = "lon_rho lat_rho benlayer ocean_time" ;
		DetBen:field = "benthic detritus, scalar, series" ;
		DetBen:_FillValue = 1.e+37f ;
	float DetF(ocean_time, s_rho, eta_rho, xi_rho) ;
		DetF:long_name = "Fast-sinking detritus concentration" ;
		DetF:units = "mg C m^-3" ;
		DetF:time = "ocean_time" ;
		DetF:grid = "grid" ;
		DetF:location = "face" ;
		DetF:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		DetF:field = "detritus, scalar, series" ;
		DetF:_FillValue = 1.e+37f ;
	double DiL ;
		DiL:long_name = "Doubling rate parameter" ;
		DiL:units = "d^-1" ;
	double DiS ;
		DiS:long_name = "Doubling rate parameter" ;
		DiS:units = "d^-1" ;
	double DpL ;
		DpL:long_name = "Doubling rate exponent" ;
		DpL:units = "degC^-1" ;
	double DpS ;
		DpS:long_name = "Doubling rate exponent" ;
		DpS:units = "degC^-1" ;
	float EupO(ocean_time, s_rho, eta_rho, xi_rho) ;
		EupO:long_name = "Offshore euphausiid concentration" ;
		EupO:units = "mg C m^-3" ;
		EupO:time = "ocean_time" ;
		EupO:grid = "grid" ;
		EupO:location = "face" ;
		EupO:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		EupO:field = "euphausiid, scalar, series" ;
		EupO:_FillValue = 1.e+37f ;
	float EupS(ocean_time, s_rho, eta_rho, xi_rho) ;
		EupS:long_name = "On-shelf euphausiid concentration" ;
		EupS:units = "mg C m^-3" ;
		EupS:time = "ocean_time" ;
		EupS:grid = "grid" ;
		EupS:location = "face" ;
		EupS:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		EupS:field = "euphausiid, scalar, series" ;
		EupS:_FillValue = 1.e+37f ;
	double FSobc_in(boundary) ;
		FSobc_in:long_name = "free-surface inflow, nudging inverse time scale" ;
		FSobc_in:units = "second-1" ;
	double FSobc_out(boundary) ;
		FSobc_out:long_name = "free-surface outflow, nudging inverse time scale" ;
		FSobc_out:units = "second-1" ;
	double Falpha ;
		Falpha:long_name = "Power-law shape barotropic filter parameter" ;
	double Fbeta ;
		Fbeta:long_name = "Power-law shape barotropic filter parameter" ;
	float Fe(ocean_time, s_rho, eta_rho, xi_rho) ;
		Fe:long_name = "Iron concentration" ;
		Fe:units = "umol Fe m^-3" ;
		Fe:time = "ocean_time" ;
		Fe:grid = "grid" ;
		Fe:location = "face" ;
		Fe:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		Fe:field = "iron conc, scalar, series" ;
		Fe:_FillValue = 1.e+37f ;
	double FeC ;
		FeC:long_name = "Fe:Carbon ratio    (2 umol Fe : mol C)" ;
		FeC:units = "umol Fe / mg C" ;
	double FeCritPL ;
		FeCritPL:long_name = "Threshold below which PhS is limited" ;
		FeCritPL:units = "umol Fe m^-3" ;
	double FeCritPS ;
		FeCritPS:long_name = "Threshold below which PhS is limited" ;
		FeCritPS:units = "umol Fe m^-3" ;
	double Feinh ;
		Feinh:long_name = "inshore isobath of transition" ;
		Feinh:units = "m" ;
	double Feinhi ;
		Feinhi:long_name = "inshore/deep" ;
		Feinhi:units = "micromol Fe m-3 or nM" ;
	double Feinlo ;
		Feinlo:long_name = "inshore/surface" ;
		Feinlo:units = "micromol Fe m-3 or nM" ;
	double Feoffh ;
		Feoffh:long_name = "offshore isobath of transition" ;
		Feoffh:units = "m" ;
	double Feoffhi ;
		Feoffhi:long_name = "offshore/deep" ;
		Feoffhi:units = "micromol Fe m-3 or nM" ;
	double Feofflo ;
		Feofflo:long_name = "offshore/surface" ;
		Feofflo:units = "micromol Fe m-3 or nM" ;
	double Fgamma ;
		Fgamma:long_name = "Power-law shape barotropic filter parameter" ;
	float Hsbl(ocean_time, eta_rho, xi_rho) ;
		Hsbl:long_name = "depth of oceanic surface boundary layer" ;
		Hsbl:units = "meter" ;
		Hsbl:time = "ocean_time" ;
		Hsbl:grid = "grid" ;
		Hsbl:location = "face" ;
		Hsbl:coordinates = "lon_rho lat_rho ocean_time" ;
		Hsbl:field = "Hsbl, scalar, series" ;
		Hsbl:_FillValue = 1.e+37f ;
	float IceNH4(ocean_time, eta_rho, xi_rho) ;
		IceNH4:long_name = "Ice ammonium concentration" ;
		IceNH4:units = "mmol N m^-3" ;
		IceNH4:time = "ocean_time" ;
		IceNH4:grid = "grid" ;
		IceNH4:location = "face" ;
		IceNH4:coordinates = "lon_rho lat_rho ocean_time" ;
		IceNH4:field = "ice ammonium conc, scalar, series" ;
		IceNH4:_FillValue = 1.e+37f ;
	float IceNO3(ocean_time, eta_rho, xi_rho) ;
		IceNO3:long_name = "Ice nitrate concentration" ;
		IceNO3:units = "mmol N m^-3" ;
		IceNO3:time = "ocean_time" ;
		IceNO3:grid = "grid" ;
		IceNO3:location = "face" ;
		IceNO3:coordinates = "lon_rho lat_rho ocean_time" ;
		IceNO3:field = "ice nitrate conc, scalar, series" ;
		IceNO3:_FillValue = 1.e+37f ;
	float IcePhL(ocean_time, eta_rho, xi_rho) ;
		IcePhL:long_name = "Ice algae concentration" ;
		IcePhL:units = "mg C m^-3" ;
		IcePhL:time = "ocean_time" ;
		IcePhL:grid = "grid" ;
		IcePhL:location = "face" ;
		IcePhL:coordinates = "lon_rho lat_rho ocean_time" ;
		IcePhL:field = "ice algae conc, scalar, series" ;
		IcePhL:_FillValue = 1.e+37f ;
	float Jel(ocean_time, s_rho, eta_rho, xi_rho) ;
		Jel:long_name = "Jellyfish concentration" ;
		Jel:units = "mg C m^-3" ;
		Jel:time = "ocean_time" ;
		Jel:grid = "grid" ;
		Jel:location = "face" ;
		Jel:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		Jel:field = "jellyfish, scalar, series" ;
		Jel:_FillValue = 1.e+37f ;
	double KI ;
		KI:long_name = "Nitrification light half-saturation constant" ;
		KI:units = "W m^-2" ;
	double KNH4Nit ;
		KNH4Nit:long_name = "Half saturation constant for nitrification" ;
		KNH4Nit:units = "mmolN/m^3" ;
	double KtBm_MZL ;
		KtBm_MZL:long_name = "temperature coefficient for respiration" ;
		KtBm_MZL:units = "1/deg C" ;
	double KtBm_PhL ;
		KtBm_PhL:long_name = "temperature coefficient for respiration" ;
		KtBm_PhL:units = "1/deg C" ;
	double KtBm_PhS ;
		KtBm_PhS:long_name = "temperature coefficient for respiration" ;
		KtBm_PhS:units = "1/deg C" ;
	double KupD ;
		KupD:long_name = "Half-saturation constant for feeding on benthic prey" ;
		KupD:units = "mg C/m^2" ;
	double KupP ;
		KupP:long_name = "Half-saturation constant for feeding on pelagic prey" ;
		KupP:units = "mg C/m^2" ;
	int Lm2CLM ;
		Lm2CLM:long_name = "2D momentum climatology processing switch" ;
		Lm2CLM:flag_values = 0, 1 ;
		Lm2CLM:flag_meanings = ".FALSE. .TRUE." ;
	int Lm3CLM ;
		Lm3CLM:long_name = "3D momentum climatology processing switch" ;
		Lm3CLM:flag_values = 0, 1 ;
		Lm3CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeM2CLM ;
		LnudgeM2CLM:long_name = "2D momentum climatology nudging activation switch" ;
		LnudgeM2CLM:flag_values = 0, 1 ;
		LnudgeM2CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeM3CLM ;
		LnudgeM3CLM:long_name = "3D momentum climatology nudging activation switch" ;
		LnudgeM3CLM:flag_values = 0, 1 ;
		LnudgeM3CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeTCLM(tracer) ;
		LnudgeTCLM:long_name = "tracer climatology nudging activation switch" ;
		LnudgeTCLM:flag_values = 0, 1 ;
		LnudgeTCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LsshCLM ;
		LsshCLM:long_name = "sea surface height climatology processing switch" ;
		LsshCLM:flag_values = 0, 1 ;
		LsshCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerCLM(tracer) ;
		LtracerCLM:long_name = "tracer climatology processing switch" ;
		LtracerCLM:flag_values = 0, 1 ;
		LtracerCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerSponge(tracer) ;
		LtracerSponge:long_name = "horizontal diffusivity sponge activation switch" ;
		LtracerSponge:flag_values = 0, 1 ;
		LtracerSponge:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerSrc(tracer) ;
		LtracerSrc:long_name = "tracer point sources and sink activation switch" ;
		LtracerSrc:flag_values = 0, 1 ;
		LtracerSrc:flag_meanings = ".FALSE. .TRUE." ;
	double LupD ;
		LupD:long_name = "Lower threshold for feeding on benthic prey" ;
		LupD:units = "mg C/m^2" ;
	double LupP ;
		LupP:long_name = "Lower threshold for feeding on pelagic prey" ;
		LupP:units = "mg C/m^2" ;
	int LuvSponge ;
		LuvSponge:long_name = "horizontal viscosity sponge activation switch" ;
		LuvSponge:flag_values = 0, 1 ;
		LuvSponge:flag_meanings = ".FALSE. .TRUE." ;
	int LuvSrc ;
		LuvSrc:long_name = "momentum point sources and sink activation switch" ;
		LuvSrc:flag_values = 0, 1 ;
		LuvSrc:flag_meanings = ".FALSE. .TRUE." ;
	int LwSrc ;
		LwSrc:long_name = "mass point sources and sink activation switch" ;
		LwSrc:flag_values = 0, 1 ;
		LwSrc:flag_meanings = ".FALSE. .TRUE." ;
	double M2nudg ;
		M2nudg:long_name = "2D momentum nudging/relaxation inverse time scale" ;
		M2nudg:units = "day-1" ;
	double M2obc_in(boundary) ;
		M2obc_in:long_name = "2D momentum inflow, nudging inverse time scale" ;
		M2obc_in:units = "second-1" ;
	double M2obc_out(boundary) ;
		M2obc_out:long_name = "2D momentum outflow, nudging inverse time scale" ;
		M2obc_out:units = "second-1" ;
	double M3nudg ;
		M3nudg:long_name = "3D momentum nudging/relaxation inverse time scale" ;
		M3nudg:units = "day-1" ;
	double M3obc_in(boundary) ;
		M3obc_in:long_name = "3D momentum inflow, nudging inverse time scale" ;
		M3obc_in:units = "second-1" ;
	double M3obc_out(boundary) ;
		M3obc_out:long_name = "3D momentum outflow, nudging inverse time scale" ;
		M3obc_out:units = "second-1" ;
	float MZL(ocean_time, s_rho, eta_rho, xi_rho) ;
		MZL:long_name = "Microzooplankton concentration" ;
		MZL:units = "mg C m^-3" ;
		MZL:time = "ocean_time" ;
		MZL:grid = "grid" ;
		MZL:location = "face" ;
		MZL:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		MZL:field = "large microzooplankton, scalar, series" ;
		MZL:_FillValue = 1.e+37f ;
	float NCaO(ocean_time, s_rho, eta_rho, xi_rho) ;
		NCaO:long_name = "Offshore large copepod concentration" ;
		NCaO:units = "mg C m^-3" ;
		NCaO:time = "ocean_time" ;
		NCaO:grid = "grid" ;
		NCaO:location = "face" ;
		NCaO:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		NCaO:field = "neocalanus, scalar, series" ;
		NCaO:_FillValue = 1.e+37f ;
	float NCaS(ocean_time, s_rho, eta_rho, xi_rho) ;
		NCaS:long_name = "On-shelf large copepod concentration" ;
		NCaS:units = "mg C m^-3" ;
		NCaS:time = "ocean_time" ;
		NCaS:grid = "grid" ;
		NCaS:location = "face" ;
		NCaS:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		NCaS:field = "neocalanus, scalar, series" ;
		NCaS:_FillValue = 1.e+37f ;
	float NH4(ocean_time, s_rho, eta_rho, xi_rho) ;
		NH4:long_name = "Ammonium concentration" ;
		NH4:units = "mmol N m^-3" ;
		NH4:time = "ocean_time" ;
		NH4:grid = "grid" ;
		NH4:location = "face" ;
		NH4:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		NH4:field = "NH4, scalar, series" ;
		NH4:_FillValue = 1.e+37f ;
	float NO3(ocean_time, s_rho, eta_rho, xi_rho) ;
		NO3:long_name = "Nitrate concentration" ;
		NO3:units = "mmol N m^-3" ;
		NO3:time = "ocean_time" ;
		NO3:grid = "grid" ;
		NO3:location = "face" ;
		NO3:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		NO3:field = "NO3, scalar, series" ;
		NO3:_FillValue = 1.e+37f ;
	double Nitr0 ;
		Nitr0:long_name = "Nitrification rate at 0C" ;
		Nitr0:units = "1/d" ;
	double PARfrac ;
		PARfrac:long_name = "Fraction of irradiance that is photosynthetically available (PAR)" ;
		PARfrac:units = "unitless" ;
	float PhL(ocean_time, s_rho, eta_rho, xi_rho) ;
		PhL:long_name = "Large phytoplankton concentration" ;
		PhL:units = "mg C m^-3" ;
		PhL:time = "ocean_time" ;
		PhL:grid = "grid" ;
		PhL:location = "face" ;
		PhL:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		PhL:field = "large phytoplankton, scalar, series" ;
		PhL:_FillValue = 1.e+37f ;
	float PhS(ocean_time, s_rho, eta_rho, xi_rho) ;
		PhS:long_name = "Small phytoplankton concentration" ;
		PhS:units = "mg C m^-3" ;
		PhS:time = "ocean_time" ;
		PhS:grid = "grid" ;
		PhS:location = "face" ;
		PhS:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		PhS:field = "small phytoplankton, scalar, series" ;
		PhS:_FillValue = 1.e+37f ;
	double Pv0 ;
		Pv0:long_name = "PON decompositon at 0 deg C" ;
		Pv0:units = "1/d" ;
	double PvT ;
		PvT:long_name = "Temperature coefficient for remineralization" ;
		PvT:units = "1/deg C" ;
	double Q10Cop ;
		Q10Cop:long_name = "Q10 for growth rate" ;
		Q10Cop:units = "unitless" ;
	double Q10CopT ;
		Q10CopT:long_name = "Temperature coefficient for Q10" ;
		Q10CopT:units = "deg. C" ;
	double Q10Eup ;
		Q10Eup:long_name = "Q10 for growth rate" ;
		Q10Eup:units = "unitless" ;
	double Q10EupT ;
		Q10EupT:long_name = "Temperature coefficient for Q10" ;
		Q10EupT:units = "deg. C" ;
	double Q10JelTe ;
		Q10JelTe:long_name = "Temperature coefficient for Q10" ;
		Q10JelTe:units = "deg. C" ;
	double Q10JelTr ;
		Q10JelTr:long_name = "reference temperature for Q10 respiration, jellyfish" ;
		Q10JelTr:units = "1/degC" ;
	double Q10Jele ;
		Q10Jele:long_name = "Q10 for growth rate" ;
		Q10Jele:units = "unitless" ;
	double Q10Jelr ;
		Q10Jelr:long_name = "Q10 for respiration rate, jellyfish" ;
		Q10Jelr:units = "degC" ;
	double Q10MZL ;
		Q10MZL:long_name = "Q10 for growth rate" ;
		Q10MZL:units = "unitless" ;
	double Q10MZLT ;
		Q10MZLT:long_name = "Temperature coefficient for Q10" ;
		Q10MZLT:units = "deg. C" ;
	double Q10NCa ;
		Q10NCa:long_name = "Q10 for growth rate" ;
		Q10NCa:units = "unitless" ;
	double Q10NCaT ;
		Q10NCaT:long_name = "Temperature coefficient for Q10" ;
		Q10NCaT:units = "deg. C" ;
	double Qres ;
		Qres:long_name = "Active metabolic rate" ;
		Qres:units = "1/d" ;
	double R0i ;
		R0i:long_name = "IcePhL respiration rate" ;
		R0i:units = "1/d" ;
	double RiseEnd ;
		RiseEnd:long_name = "Date NCaO stop moving upward" ;
		RiseEnd:units = "Day of Year" ;
	double RiseEndCM ;
		RiseEndCM:long_name = "Date NCaS stop moving upward" ;
		RiseEndCM:units = "Day of Year" ;
	double RiseStart ;
		RiseStart:long_name = "Date NCaO begin to move upward" ;
		RiseStart:units = "Day of Year" ;
	double RiseStartCM ;
		RiseStartCM:long_name = "Date NCaS begin to move upward" ;
		RiseStartCM:units = "Day of Year" ;
	double Rres ;
		Rres:long_name = "Basal metabolism rate" ;
		Rres:units = "1/d" ;
	double Rup ;
		Rup:long_name = "maximum specific ingestion rate" ;
		Rup:units = "1/d" ;
	double SinkEnd ;
		SinkEnd:long_name = "Date NCaO stop moving downward" ;
		SinkEnd:units = "Day of Year" ;
	double SinkEndCM ;
		SinkEndCM:long_name = "Date NCaS stop moving downward" ;
		SinkEndCM:units = "Day of Year" ;
	double SinkStart ;
		SinkStart:long_name = "Date NCaO begin to move downward" ;
		SinkStart:units = "Day of Year" ;
	double SinkStartCM ;
		SinkStartCM:long_name = "Date NCaS begin to move downward" ;
		SinkStartCM:units = "Day of Year" ;
	double T0benr ;
		T0benr:long_name = "Reference temperature for growth/feeding rate" ;
		T0benr:units = "degC" ;
	float TIC(ocean_time, s_rho, eta_rho, xi_rho) ;
		TIC:long_name = "total inorganic carbon" ;
		TIC:units = "mmol C m^-3" ;
		TIC:time = "ocean_time" ;
		TIC:grid = "grid" ;
		TIC:location = "face" ;
		TIC:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		TIC:field = "TIC, scalar, series" ;
		TIC:_FillValue = 1.e+37f ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double TmaxMZL ;
		TmaxMZL:long_name = "reference temperature for respiration" ;
		TmaxMZL:units = "degC" ;
	double TmaxPhL ;
		TmaxPhL:long_name = "reference temperature for respiration" ;
		TmaxPhL:units = "degC" ;
	double TmaxPhS ;
		TmaxPhS:long_name = "reference temperature for respiration" ;
		TmaxPhS:units = "degC" ;
	double Tnudg(tracer) ;
		Tnudg:long_name = "Tracers nudging/relaxation inverse time scale" ;
		Tnudg:units = "day-1" ;
	double Tnudg_SSS ;
		Tnudg_SSS:long_name = "SSS nudging/relaxation inverse time scale" ;
		Tnudg_SSS:units = "day-1" ;
	double Tobc_in(boundary, tracer) ;
		Tobc_in:long_name = "tracers inflow, nudging inverse time scale" ;
		Tobc_in:units = "second-1" ;
	double Tobc_out(boundary, tracer) ;
		Tobc_out:long_name = "tracers outflow, nudging inverse time scale" ;
		Tobc_out:units = "second-1" ;
	double ToptNtr ;
		ToptNtr:long_name = "Optimal temperature for nitrification" ;
		ToptNtr:units = "degC" ;
	double TrefC ;
		TrefC:long_name = "reference temperature for respiration" ;
		TrefC:units = "degC" ;
	double TrefE ;
		TrefE:long_name = "reference temperature for respiration" ;
		TrefE:units = "degC" ;
	double TrefN ;
		TrefN:long_name = "reference temperature for respiration" ;
		TrefN:units = "degC" ;
	int Vstretching ;
		Vstretching:long_name = "vertical terrain-following stretching function" ;
	int Vtransform ;
		Vtransform:long_name = "vertical terrain-following transformation equation" ;
	double Znudg ;
		Znudg:long_name = "free-surface nudging/relaxation inverse time scale" ;
		Znudg:units = "day-1" ;
	double Zob ;
		Zob:long_name = "bottom roughness" ;
		Zob:units = "meter" ;
	double Zos ;
		Zos:long_name = "surface roughness" ;
		Zos:units = "meter" ;
	float ageice(ocean_time, eta_rho, xi_rho) ;
		ageice:long_name = "age of the ice" ;
		ageice:units = "sec" ;
		ageice:time = "ocean_time" ;
		ageice:grid = "grid" ;
		ageice:location = "face" ;
		ageice:coordinates = "lon_rho lat_rho ocean_time" ;
		ageice:field = "ice age, scalar, series" ;
		ageice:_FillValue = 1.e+37f ;
	float aice(ocean_time, eta_rho, xi_rho) ;
		aice:long_name = "fraction of cell covered by ice" ;
		aice:time = "ocean_time" ;
		aice:grid = "grid" ;
		aice:location = "face" ;
		aice:coordinates = "lon_rho lat_rho ocean_time" ;
		aice:field = "ice concentration, scalar, series" ;
		aice:_FillValue = 1.e+37f ;
	double aidz ;
		aidz:long_name = "Ice thickness" ;
		aidz:units = "m" ;
	float alkalinity(ocean_time, s_rho, eta_rho, xi_rho) ;
		alkalinity:long_name = "total alkalinity" ;
		alkalinity:units = "mmol C m^-3" ;
		alkalinity:time = "ocean_time" ;
		alkalinity:grid = "grid" ;
		alkalinity:location = "face" ;
		alkalinity:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		alkalinity:field = "TAlk, scalar, series" ;
		alkalinity:_FillValue = 1.e+37f ;
	double alphaIb ;
		alphaIb:long_name = "IcePhL Chl-a specific attenuation coefficient" ;
		alphaIb:units = "W^-1 m^-2" ;
	double alphaPhL ;
		alphaPhL:long_name = "photosynthetic efficiency" ;
		alphaPhL:units = "mg C m^2 (mg Chl-a)^-1 (E^-1)" ;
	double alphaPhS ;
		alphaPhS:long_name = "photosynthetic efficiency" ;
		alphaPhS:units = "mg C m^2 (mg Chl-a)^-1 (E^-1)" ;
	double annit ;
		annit:long_name = "IcePhL nitrification factor" ;
		annit:units = "1/d" ;
	double betaI ;
		betaI:long_name = "IcePhL photosynthetic efficiency" ;
		betaI:units = "W^-1 m^-2" ;
	double ccr ;
		ccr:long_name = "Carbon:Chlorophyll ratio, small phyto" ;
		ccr:units = "mg C / mg Chl-a" ;
	double ccrPhL ;
		ccrPhL:long_name = "Carbon:Chlorophyll ratio, large phyto" ;
		ccrPhL:units = "mg C / mg Chl-a" ;
	float chu_iw(ocean_time, eta_rho, xi_rho) ;
		chu_iw:long_name = "ice-water momentum transfer coefficient" ;
		chu_iw:units = "meter second-1" ;
		chu_iw:time = "ocean_time" ;
		chu_iw:grid = "grid" ;
		chu_iw:location = "face" ;
		chu_iw:coordinates = "lon_rho lat_rho ocean_time" ;
		chu_iw:field = "transfer coefficient, scalar, series" ;
		chu_iw:_FillValue = 1.e+37f ;
	double dstart ;
		dstart:long_name = "time stamp assigned to model initilization" ;
		dstart:units = "days since 1900-01-01 00:00:00" ;
		dstart:calendar = "proleptic_gregorian" ;
	double dt ;
		dt:long_name = "size of long time-steps" ;
		dt:units = "second" ;
	double dtfast ;
		dtfast:long_name = "size of short time-steps" ;
		dtfast:units = "second" ;
	double eCop ;
		eCop:long_name = "maximum specific ingestion rate" ;
		eCop:units = "mg C/mg C/d" ;
	double eEup ;
		eEup:long_name = "maximum specific ingestion rate" ;
		eEup:units = "mg C/mg C/d" ;
	double eJel ;
		eJel:long_name = "maximum specific ingestion rate" ;
		eJel:units = "mg C/mg C/d" ;
	double eMZL ;
		eMZL:long_name = "maximum specific ingestion rate" ;
		eMZL:units = "mg C/mg C/d" ;
	double eNCa ;
		eNCa:long_name = "maximum specific ingestion rate" ;
		eNCa:units = "mg C/mg C/d" ;
	double eex ;
		eex:long_name = "fraction of living food excreted (1 - growth efficiency)" ;
	double eexD ;
		eexD:long_name = "fraction of detrital food excreted" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	double fCop ;
		fCop:long_name = "Half-saturation constant for grazing" ;
		fCop:units = "mg C/m3" ;
	double fEup ;
		fEup:long_name = "Half-saturation constant for grazing" ;
		fEup:units = "mg C/m3" ;
	double fJel ;
		fJel:long_name = "Half-saturation constant for grazing" ;
		fJel:units = "mg C/m3" ;
	double fMZL ;
		fMZL:long_name = "Half-saturation constant for grazing" ;
		fMZL:units = "mg C/m3" ;
	double fNCa ;
		fNCa:long_name = "Half-saturation constant for grazing" ;
		fNCa:units = "mg C/m3" ;
	double fpCopEup ;
		fpCopEup:long_name = "Cop->Eup  Feeding preference" ;
	double fpCopJel ;
		fpCopJel:long_name = "Cop->Jel  Feeding preference" ;
	double fpDetEup ;
		fpDetEup:long_name = "Det->Eup  Feeding preference" ;
	double fpDetEupO ;
		fpDetEupO:long_name = "Det->EupO Feeding preference" ;
	double fpEupJel ;
		fpEupJel:long_name = "Eup->Jel  Feeding preference" ;
	double fpMZLCop ;
		fpMZLCop:long_name = "MZL->Cop  Feeding preference" ;
	double fpMZLEup ;
		fpMZLEup:long_name = "MZL->Eup  Feeding preference" ;
	double fpMZLNCa ;
		fpMZLNCa:long_name = "MZL->NCa  Feeding preference" ;
	double fpNCaJel ;
		fpNCaJel:long_name = "NCa->Jel  Feeding preference" ;
	double fpPhLCop ;
		fpPhLCop:long_name = "PhL->Cop  Feeding preference" ;
	double fpPhLEup ;
		fpPhLEup:long_name = "PhL->Eup  Feeding preference" ;
	double fpPhLMZL ;
		fpPhLMZL:long_name = "PhL->MZL  Feeding preference" ;
	double fpPhLNCa ;
		fpPhLNCa:long_name = "PhL->NCa  Feeding preference" ;
	double fpPhSCop ;
		fpPhSCop:long_name = "PhS->Cop  Feeding preference" ;
	double fpPhSEup ;
		fpPhSEup:long_name = "PhS->Eup  Feeding preference" ;
	double fpPhSMZL ;
		fpPhSMZL:long_name = "PhS->MZL  Feeding preference" ;
	double fpPhSNCa ;
		fpPhSNCa:long_name = "PhS->NCa  Feeding preference" ;
	double gamma2 ;
		gamma2:long_name = "slipperiness parameter" ;
	double gammaCop ;
		gammaCop:long_name = "Growth efficiency" ;
	double gammaEup ;
		gammaEup:long_name = "Growth efficiency" ;
	double gammaJel ;
		gammaJel:long_name = "Growth efficiency" ;
	double gammaMZL ;
		gammaMZL:long_name = "Growth efficiency" ;
	double gammaNCa ;
		gammaNCa:long_name = "Growth efficiency" ;
	int grid ;
		grid:cf_role = "grid_topology" ;
		grid:topology_dimension = 2 ;
		grid:node_dimensions = "xi_psi eta_psi" ;
		grid:face_dimensions = "xi_rho: xi_psi (padding: both) eta_rho: eta_psi (padding: both)" ;
		grid:edge1_dimensions = "xi_u: xi_psi eta_u: eta_psi (padding: both)" ;
		grid:edge2_dimensions = "xi_v: xi_psi (padding: both) eta_v: eta_psi" ;
		grid:node_coordinates = "lon_psi lat_psi" ;
		grid:face_coordinates = "lon_rho lat_rho" ;
		grid:edge1_coordinates = "lon_u lat_u" ;
		grid:edge2_coordinates = "lon_v lat_v" ;
		grid:vertical_dimensions = "s_rho: s_w (padding: none)" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	float hice(ocean_time, eta_rho, xi_rho) ;
		hice:long_name = "average ice thickness in cell" ;
		hice:units = "meter" ;
		hice:time = "ocean_time" ;
		hice:grid = "grid" ;
		hice:location = "face" ;
		hice:coordinates = "lon_rho lat_rho ocean_time" ;
		hice:field = "ice thickness, scalar, series" ;
		hice:_FillValue = 1.e+37f ;
	double inhib ;
		inhib:long_name = "IcePhL NH4 inhibition on NO3 uptake" ;
		inhib:units = "m^3/mmol N" ;
	double k1PhL ;
		k1PhL:long_name = "Half-saturation constant for NO3 limitation" ;
	double k1PhS ;
		k1PhS:long_name = "Half-saturation constant for NO3 limitation" ;
	double k2PhL ;
		k2PhL:long_name = "Half-saturation constant for NH4 limitation" ;
	double k2PhS ;
		k2PhS:long_name = "Half-saturation constant for NH4 limitation" ;
	double k_chlA ;
		k_chlA:long_name = "Chlorophyll attenuation coefficient, factor" ;
		k_chlA:units = "m^-1" ;
	double k_chlB ;
		k_chlB:long_name = "Chlorophyll attenuation coefficient, exponent" ;
		k_chlB:units = "unitless" ;
	double k_chlC ;
		k_chlC:long_name = "Other material (CDOM,sediment,etc.) attenuation coefficient" ;
		k_chlC:units = "m^-1" ;
	double k_ext ;
		k_ext:long_name = "Clear-water attenuation coefficient" ;
		k_ext:units = "m^-1" ;
	double k_sed1 ;
		k_sed1:long_name = "Depth-based attenuation coefficient, factor" ;
		k_sed1:units = "m^-1" ;
	double k_sed2 ;
		k_sed2:long_name = "Depth-based attenuation coefficient, exponent" ;
		k_sed2:units = "unitless" ;
	double kfePhL ;
		kfePhL:long_name = "Half-saturation constant for Fe" ;
		kfePhL:units = "umol m^-3" ;
	double kfePhS ;
		kfePhS:long_name = "Half-saturation constant for Fe" ;
		kfePhS:units = "umol m^-3" ;
	double ksnut1 ;
		ksnut1:long_name = "IcePhL half-saturation constant for NO3" ;
		ksnut1:units = "mmolN/m^3" ;
	double ksnut2 ;
		ksnut2:long_name = "IcePhL half-saturation constant for NH4" ;
		ksnut2:units = "mmolN/m^3" ;
	double ktbmC ;
		ktbmC:long_name = "temperature coefficient for respiration" ;
		ktbmC:units = "1/deg C" ;
	double ktbmE ;
		ktbmE:long_name = "temperature coefficient for respiration" ;
		ktbmE:units = "1/deg C" ;
	double ktbmN ;
		ktbmN:long_name = "temperature coefficient for respiration" ;
		ktbmN:units = "1/deg C" ;
	double ktntr ;
		ktntr:long_name = "Temperature coefficient for nitrification" ;
		ktntr:units = "1/deg C" ;
	double mMZL ;
		mMZL:long_name = "daily linear mortality rate" ;
		mMZL:units = "1/d" ;
	double mPhL ;
		mPhL:long_name = "daily linear mortality rate (senescence)" ;
		mPhL:units = "1/d" ;
	double mPhS ;
		mPhS:long_name = "daily linear mortality rate (senescence)" ;
		mPhS:units = "1/d" ;
	double mpredCop ;
		mpredCop:long_name = "Daily mortality for Copepods" ;
		mpredCop:units = "1/d/mgC" ;
	double mpredEup ;
		mpredEup:long_name = "Daily mortality for Euphausiids" ;
		mpredEup:units = "1/d/mgC" ;
	double mpredJel ;
		mpredJel:long_name = "Daily mortality for Large Microzoo." ;
		mpredJel:units = "1/d/mgC" ;
	double mpredMZL ;
		mpredMZL:long_name = "Daily mortality for Large Microzoo." ;
		mpredMZL:units = "1/d/mgC" ;
	double mpredNCa ;
		mpredNCa:long_name = "Daily mortality for Neocalanus" ;
		mpredNCa:units = "1/d/mgC" ;
	double mu0 ;
		mu0:long_name = "IcePhL maximum growth rate at 0 deg C" ;
		mu0:units = "1/d" ;
	int nAVG ;
		nAVG:long_name = "number of time-steps between time-averaged records" ;
	int nDIA ;
		nDIA:long_name = "number of time-steps between diagnostic records" ;
	int nHIS ;
		nHIS:long_name = "number of time-steps between history records" ;
	int nRST ;
		nRST:long_name = "number of time-steps between restart records" ;
		nRST:cycle = "only latest two records are maintained" ;
	int nSTA ;
		nSTA:long_name = "number of time-steps between stations records" ;
	int ndefAVG ;
		ndefAVG:long_name = "number of time-steps between the creation of average files" ;
	int ndefDIA ;
		ndefDIA:long_name = "number of time-steps between the creation of diagnostic files" ;
	int ndefHIS ;
		ndefHIS:long_name = "number of time-steps between the creation of history files" ;
	int ndtfast ;
		ndtfast:long_name = "number of short time-steps" ;
	double nl_tnu2(tracer) ;
		nl_tnu2:long_name = "nonlinear model Laplacian mixing coefficient for tracers" ;
		nl_tnu2:units = "meter2 second-1" ;
	double nl_visc2 ;
		nl_visc2:long_name = "nonlinear model Laplacian mixing coefficient for momentum" ;
		nl_visc2:units = "meter2 second-1" ;
	int ntimes ;
		ntimes:long_name = "number of long time-steps" ;
	int ntsAVG ;
		ntsAVG:long_name = "starting time-step for accumulation of time-averaged fields" ;
	int ntsDIA ;
		ntsDIA:long_name = "starting time-step for accumulation of diagnostic fields" ;
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 1900-01-01 00:00:00" ;
		ocean_time:calendar = "proleptic_gregorian" ;
		ocean_time:field = "time, scalar, series" ;
	float oxygen(ocean_time, s_rho, eta_rho, xi_rho) ;
		oxygen:long_name = "dissolved oxygen concentration" ;
		oxygen:units = "mmol O m^-3" ;
		oxygen:time = "ocean_time" ;
		oxygen:grid = "grid" ;
		oxygen:location = "face" ;
		oxygen:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		oxygen:field = "Oxygen, scalar, series" ;
		oxygen:_FillValue = 1.e+37f ;
	double prefD ;
		prefD:long_name = "DetBen->Ben feeding preference" ;
	double prefPL ;
		prefPL:long_name = "PhL->Ben feeding preference" ;
	double prefPS ;
		prefPS:long_name = "PhS->Ben feeding preference" ;
	double q10r ;
		q10r:long_name = "Q10 for growth/feeding and mortality rate" ;
		q10r:units = "unitless" ;
	double rdrg ;
		rdrg:long_name = "linear drag coefficient" ;
		rdrg:units = "meter second-1" ;
	double rdrg2 ;
		rdrg2:long_name = "quadratic drag coefficient" ;
	double respCop ;
		respCop:long_name = "Specific respiration rate" ;
		respCop:units = "d^-1" ;
	double respEup ;
		respEup:long_name = "Specific respiration rate" ;
		respEup:units = "d^-1" ;
	double respJel ;
		respJel:long_name = "Specific respiration rate" ;
		respJel:units = "d^-1" ;
	double respMZL ;
		respMZL:long_name = "Specific respiration rate" ;
		respMZL:units = "d^-1" ;
	double respNCa ;
		respNCa:long_name = "Specific respiration rate" ;
		respNCa:units = "d^-1" ;
	double respPhL ;
		respPhL:long_name = "Specific respiration rate" ;
		respPhL:units = "d^-1" ;
	double respPhS ;
		respPhS:long_name = "Specific respiration rate" ;
		respPhS:units = "d^-1" ;
	double rg ;
		rg:long_name = "IcePhL temperature coefficient for mortality" ;
		rg:units = "1/deg C" ;
	double rg0 ;
		rg0:long_name = "IcePhL mortality rate at 0 deg C" ;
		rg0:units = "1/d" ;
	float rho(ocean_time, s_rho, eta_rho, xi_rho) ;
		rho:long_name = "density anomaly" ;
		rho:units = "kilogram meter-3" ;
		rho:time = "ocean_time" ;
		rho:grid = "grid" ;
		rho:location = "face" ;
		rho:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		rho:field = "density, scalar, series" ;
		rho:_FillValue = 1.e+37f ;
	double rho0 ;
		rho0:long_name = "mean density used in Boussinesq approximation" ;
		rho0:units = "kilogram meter-3" ;
	double rmort ;
		rmort:long_name = "linear mortality rate" ;
		rmort:units = "1/d" ;
	float s0mk(ocean_time, eta_rho, xi_rho) ;
		s0mk:long_name = "salinity of molecular sub-layer under ice" ;
		s0mk:time = "ocean_time" ;
		s0mk:grid = "grid" ;
		s0mk:location = "face" ;
		s0mk:coordinates = "lon_rho lat_rho ocean_time" ;
		s0mk:field = "salinity, scalar, series" ;
		s0mk:_FillValue = 1.e+37f ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
		s_rho:positive = "up" ;
		s_rho:standard_name = "ocean_s_coordinate_g1" ;
		s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
		s_rho:field = "s_rho, scalar" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
		s_w:positive = "up" ;
		s_w:standard_name = "ocean_s_coordinate_g1" ;
		s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
		s_w:field = "s_w, scalar" ;
	float salt(ocean_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:time = "ocean_time" ;
		salt:grid = "grid" ;
		salt:location = "face" ;
		salt:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		salt:field = "salinity, scalar, series" ;
		salt:_FillValue = 1.e+37f ;
	float sig11(ocean_time, eta_rho, xi_rho) ;
		sig11:long_name = "internal ice stress 11 component" ;
		sig11:units = "Newton meter-1" ;
		sig11:time = "ocean_time" ;
		sig11:grid = "grid" ;
		sig11:location = "face" ;
		sig11:coordinates = "lon_rho lat_rho ocean_time" ;
		sig11:field = "ice stress 11, scalar, series" ;
		sig11:_FillValue = 1.e+37f ;
	float sig12(ocean_time, eta_rho, xi_rho) ;
		sig12:long_name = "internal ice stress 12 component" ;
		sig12:units = "Newton meter-1" ;
		sig12:time = "ocean_time" ;
		sig12:grid = "grid" ;
		sig12:location = "face" ;
		sig12:coordinates = "lon_rho lat_rho ocean_time" ;
		sig12:field = "ice stress 12, scalar, series" ;
		sig12:_FillValue = 1.e+37f ;
	float sig22(ocean_time, eta_rho, xi_rho) ;
		sig22:long_name = "internal ice stress 22 component" ;
		sig22:units = "Newton meter-1" ;
		sig22:time = "ocean_time" ;
		sig22:grid = "grid" ;
		sig22:location = "face" ;
		sig22:coordinates = "lon_rho lat_rho ocean_time" ;
		sig22:field = "ice stress 22, scalar, series" ;
		sig22:_FillValue = 1.e+37f ;
	float snow_thick(ocean_time, eta_rho, xi_rho) ;
		snow_thick:long_name = "thickness of snow cover" ;
		snow_thick:units = "meter" ;
		snow_thick:time = "ocean_time" ;
		snow_thick:grid = "grid" ;
		snow_thick:location = "face" ;
		snow_thick:coordinates = "lon_rho lat_rho ocean_time" ;
		snow_thick:field = "snow thickness, scalar, series" ;
		snow_thick:_FillValue = 1.e+37f ;
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = 0, 1 ;
		spherical:flag_meanings = "Cartesian spherical" ;
	float t0mk(ocean_time, eta_rho, xi_rho) ;
		t0mk:long_name = "temperature of molecular sub-layer under ice" ;
		t0mk:units = "degrees Celsius" ;
		t0mk:time = "ocean_time" ;
		t0mk:grid = "grid" ;
		t0mk:location = "face" ;
		t0mk:coordinates = "lon_rho lat_rho ocean_time" ;
		t0mk:field = "temperature, scalar, series" ;
		t0mk:_FillValue = 1.e+37f ;
	double tI0 ;
		tI0:long_name = "Nitrification light threshold" ;
		tI0:units = "W m^-2" ;
	float tau_iw(ocean_time, eta_rho, xi_rho) ;
		tau_iw:long_name = "ice-water friction velocity" ;
		tau_iw:units = "meter second-1" ;
		tau_iw:time = "ocean_time" ;
		tau_iw:grid = "grid" ;
		tau_iw:location = "face" ;
		tau_iw:coordinates = "lon_rho lat_rho ocean_time" ;
		tau_iw:field = "friction velocity, scalar, series" ;
		tau_iw:_FillValue = 1.e+37f ;
	float temp(ocean_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:time = "ocean_time" ;
		temp:grid = "grid" ;
		temp:location = "face" ;
		temp:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		temp:field = "temperature, scalar, series" ;
		temp:_FillValue = 1.e+37f ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	float ti(ocean_time, eta_rho, xi_rho) ;
		ti:long_name = "interior ice temperature" ;
		ti:units = "degrees Celcius" ;
		ti:time = "ocean_time" ;
		ti:grid = "grid" ;
		ti:location = "face" ;
		ti:coordinates = "lon_rho lat_rho ocean_time" ;
		ti:field = "interior temperature, scalar, series" ;
		ti:_FillValue = 1.e+37f ;
	float tisrf(ocean_time, eta_rho, xi_rho) ;
		tisrf:long_name = "temperature of ice surface" ;
		tisrf:units = "degrees Celcius" ;
		tisrf:time = "ocean_time" ;
		tisrf:grid = "grid" ;
		tisrf:location = "face" ;
		tisrf:coordinates = "lon_rho lat_rho ocean_time" ;
		tisrf:field = "surface temperature, scalar, series" ;
		tisrf:_FillValue = 1.e+37f ;
	float u(ocean_time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:time = "ocean_time" ;
		u:grid = "grid" ;
		u:location = "edge1" ;
		u:coordinates = "lon_u lat_u s_rho ocean_time" ;
		u:field = "u-velocity, scalar, series" ;
		u:_FillValue = 1.e+37f ;
	float ubar(ocean_time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:time = "ocean_time" ;
		ubar:grid = "grid" ;
		ubar:location = "edge1" ;
		ubar:coordinates = "lon_u lat_u ocean_time" ;
		ubar:field = "ubar-velocity, scalar, series" ;
		ubar:_FillValue = 1.e+37f ;
	float uice(ocean_time, eta_u, xi_u) ;
		uice:long_name = "u-component of ice velocity" ;
		uice:units = "meter second-1" ;
		uice:time = "ocean_time" ;
		uice:grid = "grid" ;
		uice:location = "edge1" ;
		uice:coordinates = "lon_u lat_u ocean_time" ;
		uice:field = "u-component of ice velocity, scalar, series" ;
		uice:_FillValue = 1.e+37f ;
	float v(ocean_time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:time = "ocean_time" ;
		v:grid = "grid" ;
		v:location = "edge2" ;
		v:coordinates = "lon_v lat_v s_rho ocean_time" ;
		v:field = "v-velocity, scalar, series" ;
		v:_FillValue = 1.e+37f ;
	float vbar(ocean_time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:time = "ocean_time" ;
		vbar:grid = "grid" ;
		vbar:location = "edge2" ;
		vbar:coordinates = "lon_v lat_v ocean_time" ;
		vbar:field = "vbar-velocity, scalar, series" ;
		vbar:_FillValue = 1.e+37f ;
	float vice(ocean_time, eta_v, xi_v) ;
		vice:long_name = "v-component of ice velocity" ;
		vice:units = "meter second-1" ;
		vice:time = "ocean_time" ;
		vice:grid = "grid" ;
		vice:location = "edge2" ;
		vice:coordinates = "lon_v lat_v ocean_time" ;
		vice:field = "v-component of ice velocity, scalar, series" ;
		vice:_FillValue = 1.e+37f ;
	double wDet ;
		wDet:long_name = "Sinking rate for Detritus" ;
		wDet:units = "m/d" ;
	double wDetF ;
		wDetF:long_name = "Sinking rate for Detritus" ;
		wDetF:units = "m/d" ;
	double wNCrise ;
		wNCrise:long_name = "upward velocity , tuned not data" ;
		wNCrise:units = "m/day" ;
	double wNCsink ;
		wNCsink:long_name = "downward velocity , tuned not data" ;
		wNCsink:units = "m/day" ;
	double wPhL ;
		wPhL:long_name = "Sinking rate for Large Phytoplankton" ;
		wPhL:units = "m/d" ;
	double wPhS ;
		wPhS:long_name = "Sinking rate for Small Phytoplankton" ;
		wPhS:units = "m/d" ;
	double xi ;
		xi:long_name = "Nitrogen:Carbon ratio" ;
		xi:units = "mmol N / mg C" ;
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	float zeta(ocean_time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:units = "meter" ;
		zeta:time = "ocean_time" ;
		zeta:grid = "grid" ;
		zeta:location = "face" ;
		zeta:coordinates = "lon_rho lat_rho ocean_time" ;
		zeta:field = "free-surface, scalar, series" ;
		zeta:_FillValue = 1.e+37f ;

// global attributes:
		:file = "bgcmip_bestnpz/Out/bgcmip_bestnpz_23_rst.nc" ;
		:format = "netCDF-3 64bit offset file" ;
		:Conventions = "CF-1.4, SGRID-0.3" ;
		:type = "ROMS/TOMS restart file" ;
		:title = "Bering Sea 10km Grid" ;
		:var_info = "../bering-Apps/Apps/Bering_BGC_variants/varinfo_bestnpz_scaledbry.dat" ;
		:rst_file = "bgcmip_bestnpz/Out/bgcmip_bestnpz_23_rst.nc" ;
		:his_base = "bgcmip_bestnpz/Out/bgcmip_bestnpz_his" ;
		:avg_base = "bgcmip_bestnpz/Out/bgcmip_bestnpz_avg" ;
		:dia_base = "bgcmip_bestnpz/Out/bgcmip_bestnpz_dia" ;
		:sta_file = "bgcmip_bestnpz/Out/bgcmip_bestnpz_23_sta.nc" ;
		:grd_file = "../../ROMS_Datasets/grids/AlaskaGrids_Bering10K.nc" ;
		:ini_file = "bgcmip_bestnpz/Out/bgcmip_bestnpz_22_rst.nc" ;
		:tide_file = "../../ROMS_Datasets/OTPS/tides_OTPS_Bering10K.nc" ;
		:frc_file_01 = "../../ROMS_Datasets/BarrowCO2/atmo_co2_barrow_1970_2020.nc" ;
		:frc_file_02 = "../../ROMS_Datasets/Iron/ESM4_Bering10K_iron_dust_clim.nc" ;
		:frc_file_03 = "../../ROMS_Datasets/salinity/sss.clim.nc" ;
		:frc_file_04 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Pair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Pair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Pair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Pair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Pair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Pair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Pair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Pair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Pair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Pair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Pair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Pair-2020.nc" ;
		:frc_file_05 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Qair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Qair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Qair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Qair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Qair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Qair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Qair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Qair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Qair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Qair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Qair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Qair-2020.nc" ;
		:frc_file_06 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Tair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Tair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Tair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Tair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Tair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Tair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Tair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Tair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Tair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Tair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Tair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Tair-2020.nc" ;
		:frc_file_07 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Uwind-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Uwind-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Uwind-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Uwind-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Uwind-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Uwind-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Uwind-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Uwind-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Uwind-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Uwind-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Uwind-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Uwind-2020.nc" ;
		:frc_file_08 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Vwind-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Vwind-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Vwind-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Vwind-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Vwind-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Vwind-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Vwind-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Vwind-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Vwind-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Vwind-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Vwind-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Vwind-2020.nc" ;
		:frc_file_09 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-rain-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-rain-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-rain-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-rain-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-rain-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-rain-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-rain-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-rain-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-rain-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-rain-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-rain-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-rain-2020.nc" ;
		:frc_file_10 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-swrad-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-swrad-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-swrad-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-swrad-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-swrad-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-swrad-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-swrad-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-swrad-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-swrad-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-swrad-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-swrad-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-swrad-2020.nc" ;
		:frc_file_11 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-lwrad-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-lwrad-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-lwrad-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-lwrad-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-lwrad-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-lwrad-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-lwrad-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-lwrad-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-lwrad-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-lwrad-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-lwrad-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-lwrad-2020.nc" ;
		:frc_file_12 = "../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2009.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2010.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2011.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2012.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2013.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2014.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2015.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2016.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2017.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2018.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2019.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2020.nc" ;
		:frc_file_13 = "../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2009.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2010.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2011.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2012.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2013.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2014.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2015.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2016.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2017.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2018.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2019.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2020.nc" ;
		:bry_file_01 = "../../ROMS_Datasets/WOA2018/WOA2018_Bering10K_N30_brybgc.nc" ;
		:bry_file_02 = "../../ROMS_Datasets/CFS/2009/CFS-ocean-Bering10K-N30-bryocn-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-ocean-Bering10K-N30-bryocn-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-ocean-Bering10K-N30-bryocn-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-ocean-Bering10K-N30-bryocn-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-ocean-Bering10K-N30-bryocn-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-ocean-Bering10K-N30-bryocn-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-ocean-Bering10K-N30-bryocn-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-ocean-Bering10K-N30-bryocn-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-ocean-Bering10K-N30-bryocn-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-ocean-Bering10K-N30-bryocn-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-ocean-Bering10K-N30-bryocn-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-ocean-Bering10K-N30-bryocn-2020.nc" ;
		:bry_file_03 = "../../ROMS_Datasets/CFS/2009/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2020.nc" ;
		:script_file = "bgcmip_bestnpz/In/bgcmip_bestnpz_23_ocean.in" ;
		:bpar_file = "bgcmip_bestnpz/In/bgcmip_bestnpz_bpar.in" ;
		:spos_file = "bgcmip_bestnpz/In/bgcmip_bestnpz_spos.in" ;
		:NLM_TADV = "\n",
			"ADVECTION:   HORIZONTAL   VERTICAL     \n",
			"temp:        Centered4    Centered4    \n",
			"salt:        Centered4    Centered4    \n",
			"NO3:         HSIMT        HSIMT        \n",
			"NH4:         HSIMT        HSIMT        \n",
			"PhS:         HSIMT        HSIMT        \n",
			"PhL:         HSIMT        HSIMT        \n",
			"MZL:         HSIMT        HSIMT        \n",
			"Cop:         HSIMT        HSIMT        \n",
			"NCaS:        HSIMT        HSIMT        \n",
			"EupS:        HSIMT        HSIMT        \n",
			"NCaO:        HSIMT        HSIMT        \n",
			"EupO:        HSIMT        HSIMT        \n",
			"Det:         HSIMT        HSIMT        \n",
			"DetF:        HSIMT        HSIMT        \n",
			"Jel:         HSIMT        HSIMT        \n",
			"Fe:          HSIMT        HSIMT        \n",
			"TIC:         HSIMT        HSIMT        \n",
			"alkalinity:  HSIMT        HSIMT        \n",
			"oxygen:      HSIMT        HSIMT" ;
		:NLM_LBC = "\n",
			"EDGE:        WEST   SOUTH  EAST   NORTH  \n",
			"zeta:        Che    Che    Clo    Clo    \n",
			"ubar:        Fla    Fla    Clo    Clo    \n",
			"vbar:        Fla    Fla    Clo    Clo    \n",
			"u:           RadNud RadNud Clo    Clo    \n",
			"v:           RadNud RadNud Clo    Clo    \n",
			"temp:        RadNud RadNud Clo    Clo    \n",
			"salt:        RadNud RadNud Clo    Clo    \n",
			"NO3:         RadNud RadNud Clo    Clo    \n",
			"NH4:         RadNud RadNud Clo    Clo    \n",
			"PhS:         RadNud RadNud Clo    Clo    \n",
			"PhL:         RadNud RadNud Clo    Clo    \n",
			"MZL:         RadNud RadNud Clo    Clo    \n",
			"Cop:         RadNud RadNud Clo    Clo    \n",
			"NCaS:        RadNud RadNud Clo    Clo    \n",
			"EupS:        RadNud RadNud Clo    Clo    \n",
			"NCaO:        RadNud RadNud Clo    Clo    \n",
			"EupO:        RadNud RadNud Clo    Clo    \n",
			"Det:         RadNud RadNud Clo    Clo    \n",
			"DetF:        RadNud RadNud Clo    Clo    \n",
			"Jel:         RadNud RadNud Clo    Clo    \n",
			"Fe:          RadNud RadNud Clo    Clo    \n",
			"TIC:         RadNud RadNud Clo    Clo    \n",
			"alkalinity:  RadNud RadNud Clo    Clo    \n",
			"oxygen:      RadNud RadNud Clo    Clo    \n",
			"uice:        Gra    Gra    Clo    Clo    \n",
			"vice:        Gra    Gra    Clo    Clo    \n",
			"aice:        Clo    Clo    Clo    Clo    \n",
			"hice:        Clo    Clo    Clo    Clo    \n",
			"tisrf:       Clo    Clo    Clo    Clo    \n",
			"snow_thick:  Clo    Clo    Clo    Clo    \n",
			"sig11:       Clo    Clo    Clo    Clo    \n",
			"sig12:       Clo    Clo    Clo    Clo    \n",
			"sig22:       Clo    Clo    Clo    Clo    \n",
			"IcePhL:      Clo    Clo    Clo    Clo    \n",
			"IceNO3:      Clo    Clo    Clo    Clo    \n",
			"IceNH4:      Clo    Clo    Clo    Clo" ;
		:git_url = "git@github.com:beringnpz/roms.git" ;
		:git_rev = "cobalttweaks commit 45e0c09b9385937a8121ec16b429729e0765d253" ;
		:code_dir = "/gscratch/bumblereem/kearney/roms-kate-ice" ;
		:header_dir = "/gscratch/bumblereem/kearney/BGC_hindcasts_workdir" ;
		:header_file = "bering_10k.h" ;
		:os = "Linux" ;
		:cpu = "x86_64" ;
		:compiler_system = "ifort" ;
		:compiler_command = "/gscratch/sw/intel-201703/compilers_and_libraries_2017.2.174/linux/mpi/intel64/b" ;
		:compiler_flags = "-fp-model precise -heap-arrays -ip -O3 -traceback -check uninit -ip -O3" ;
		:tiling = "007x020" ;
		:history = "Fri Sep 22 11:02:55 2023: ncks -F -d ocean_time,1,1 /gscratch/bumblereem/kearney/BGC_hindcasts_workdir/bgcmip_bestnpz/Out/bgcmip_bestnpz_23_rst.nc ../ini_hindcastloop2_BEST_NPZ.nc\n",
			"ROMS/TOMS, Version 3.9, Tuesday - June 27, 2023 - 11:54:59 AM" ;
		:ana_file = "ROMS/Functionals/ana_btflux.h, /gscratch/bumblereem/kearney/BGC_hindcasts_workdir/ana_psource.h, ROMS/Functionals/ana_srflux.h, ROMS/Functionals/ana_stflux.h, ROMS/Functionals/ana_aiobc.h, ROMS/Functionals/ana_hiobc.h, ROMS/Functionals/ana_hsnobc.h, ROMS/Functionals/ana_itobc.h" ;
		:bio_file = "ROMS/Nonlinear/Biology/bestnpz.h" ;
		:CPP_options = "BERING_10K, ADD_FSOBC, ADD_M2OBC, ALBEDO_CURVE, ANA_BPFLUX, ANA_BSFLUX, ANA_BTFLUX, ANA_PSOURCE, ANA_SPFLUX, ASSUMED_SHAPE, AVERAGES, BEST_NPZ, !BOUNDARY_ALLGATHER, BULK_FLUXES, CARBON, CARBON_FLUX, CCSM_FLUXES, COLLECT_ALLGATHER, COASTAL_ATTEN, CORE_FORCING, CURVGRID, DIAGNOSTICS_BIO, DIAGNOSTICS_TS, DIAPAUSE, DIAPAUSE, DIFF_GRID, DIURNAL_SRFLUX, DJ_GRADPS, DOUBLE_PRECISION, EMINUSP, ICE_ADVECT, ICE_BULK_FLUXES, ICE_EVP, ICE_MK, ICE_MODEL, ICE_MOMENTUM, ICE_SMOLAR, ICE_THERMO, IRON_LIMIT, LIMIT_BSTRESS, LMD_CONVEC, LMD_MIXING, LMD_NONLOCAL, LMD_RIMIX, LMD_SHAPIRO, LMD_SKPP, LONGWAVE_OUT, MASKING, MIX_GEO_TS, MIX_S_UV, MPI, NONLINEAR, NONLIN_EOS, NO_WRITE_GRID, OPTIC_MANIZZA, !OCMIP_OXYGEN_SC, OXYGEN, POT_TIDES, POWER_LAW, PROFILE, RADIATION_2D, REDUCE_ALLGATHER, RUNOFF, RST_SINGLE, SALINITY, SCORRECTION, SOLAR_SOURCE, SOLVE3D, SSH_TIDES, STATIONS, TIDES_ASTRO, TS_DIF2, UV_ADV, UV_COR, UV_U3HADVECTION, UV_SADVECTION, UV_DRAG_GRID, UV_LDRAG, UV_TIDES, UV_VIS2, UV_SMAGORINSKY, VAR_RHO_2D, VISC_GRID, VISC_3DCOEF" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
