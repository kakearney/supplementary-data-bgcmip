netcdf CFS-atmos-northPacific-Vwind-1997 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:27 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1997/roms-cfs-atmos-Vwind-1997.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1997/CFS-atmos-northPacific-Vwind-1997.nc\n",
			"Mon Sep 10 13:43:39 2018: Time overhang added\n",
			"Mon Sep 10 13:43:35 2018: ncrcat /tmp/tp22e41aee_1037_46f1_a32a_f259abe252c7.nc frc/roms-cfs-atmos-Vwind-1997.nc /tmp/tpa8d97552_bd4a_4622_b3cd_6618b29dbc28.nc /tmp/tp621b3c94_ad85_458b_94f3_1cd66c260339.nc\n",
			"Mon Sep 10 13:43:35 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-1997.nc /tmp/tp22e41aee_1037_46f1_a32a_f259abe252c7.nc\n",
			"Thu Sep  6 10:12:11 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1997_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-1997.nc\n",
			"04-Oct-2017 17:43:05: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
