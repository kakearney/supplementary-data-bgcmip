netcdf CFS-atmos-northPacific-lwrad-2013 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	lrf_time = UNLIMITED ; // (1448 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:23:21 2022: ncks -F -O -d lrf_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2013/roms-cfs-atmos-lwrad-2013.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-lwrad-2013.nc\n",
			"Mon Sep 10 13:48:31 2018: Time overhang added\n",
			"Mon Sep 10 13:48:23 2018: ncrcat /tmp/tp9419abbe_9df1_40ea_bb0f_58099677dffc.nc frc/roms-cfs-atmos-lwrad-2013.nc /tmp/tpc8d8a6cf_d953_4dc9_9db7_97c9f019f5e2.nc /tmp/tp53c7e0e6_a025_4e50_a0ae_25a63d19b35d.nc\n",
			"Mon Sep 10 13:48:22 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2013.nc /tmp/tp9419abbe_9df1_40ea_bb0f_58099677dffc.nc\n",
			"Thu Sep  6 13:03:51 2018: ncks -O -F -d lrf_time,2,1449 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2013_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2013.nc\n",
			"04-Oct-2017 18:22:48: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
