netcdf CFS-atmos-northPacific-rain-1999 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:48:02 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1999/roms-cfs-atmos-rain-1999.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1999/CFS-atmos-northPacific-rain-1999.nc\n",
			"Mon Sep 10 13:50:06 2018: Time overhang added\n",
			"Mon Sep 10 13:50:03 2018: ncrcat /tmp/tp5061aeb0_368d_4905_967a_873a121e39ea.nc frc/roms-cfs-atmos-rain-1999.nc /tmp/tp039803cc_f4f4_4f1d_a2c0_304a37617eb6.nc /tmp/tp40d6b87f_1a1c_4a40_9277_4af2768ccc85.nc\n",
			"Mon Sep 10 13:50:02 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-1999.nc /tmp/tp5061aeb0_368d_4905_967a_873a121e39ea.nc\n",
			"Thu Sep  6 10:26:47 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1999_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-1999.nc\n",
			"04-Oct-2017 17:48:47: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
