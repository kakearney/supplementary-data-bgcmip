netcdf CFS-atmos-northPacific-Qair-2006 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:52:24 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2006/roms-cfs-atmos-Qair-2006.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2006/CFS-atmos-northPacific-Qair-2006.nc\n",
			"Mon Sep 10 13:35:33 2018: Time overhang added\n",
			"Mon Sep 10 13:35:29 2018: ncrcat /tmp/tpb042406f_e237_40e3_a42b_9f08134c40ca.nc frc/roms-cfs-atmos-Qair-2006.nc /tmp/tp9663d09b_c88c_48ab_9648_1bc87e31b75a.nc /tmp/tpe4f8075a_c5d1_4c4c_9a8a_368c8a240a52.nc\n",
			"Mon Sep 10 13:35:29 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2006.nc /tmp/tpb042406f_e237_40e3_a42b_9f08134c40ca.nc\n",
			"Thu Sep  6 11:33:24 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2006.nc\n",
			"Thu Sep  6 11:32:17 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2006_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2006.nc\n",
			"04-Oct-2017 18:03:25: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
