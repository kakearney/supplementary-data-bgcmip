netcdf CFS-atmos-northPacific-Vwind-2006 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:52:44 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2006/roms-cfs-atmos-Vwind-2006.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2006/CFS-atmos-northPacific-Vwind-2006.nc\n",
			"Mon Sep 10 13:44:30 2018: Time overhang added\n",
			"Mon Sep 10 13:44:26 2018: ncrcat /tmp/tp36e507ed_9893_48c5_b83f_a4a9e9a16dd4.nc frc/roms-cfs-atmos-Vwind-2006.nc /tmp/tp82b5228f_a604_49e3_844b_3597218c3ce9.nc /tmp/tp4327f0ee_b1ad_4e86_889a_33f3ff2311cb.nc\n",
			"Mon Sep 10 13:44:26 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2006.nc /tmp/tp36e507ed_9893_48c5_b83f_a4a9e9a16dd4.nc\n",
			"Thu Sep  6 11:37:36 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2006_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2006.nc\n",
			"04-Oct-2017 18:04:32: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
