netcdf CFS-atmos-northPacific-Pair-1991 {
dimensions:
	pair_time = UNLIMITED ; // (1459 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:missing_value = -1.e+34 ;
		Pair:_FillValue = -1.e+34 ;
		Pair:time = "pair_time" ;
		Pair:coordinates = "lon lat" ;
		Pair:long_name = "atmos pressure" ;
		Pair:history = "From roms-cfs-atmos-Pair-1991" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double pair_time(pair_time) ;
		pair_time:units = "day since 1900-01-01 00:00:00" ;
		pair_time:time_origin = "01-JAN-1900 00:00:00" ;
		pair_time:axis = "T" ;
		pair_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:25:58 2022: ncks -F -O -d pair_time,2,1460 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Pair-1991.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1991/CFS-atmos-northPacific-Pair-1991.nc\n",
			"Wed Nov 20 13:58:29 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:58:25 2019: ncrcat /tmp/tp5df2af53_3841_45fb_9f89_5c2074cf5488.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Pair-1991.nc /tmp/tp9c003191_813d_4548_8425_370a117a5f4f.nc /tmp/tpbbe97454_d7c5_4e6d_96eb_4448ef20a6bb.nc\n",
			"Wed Nov 20 13:58:23 2019: ncks -F -d pair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Pair-1991.nc /tmp/tp5df2af53_3841_45fb_9f89_5c2074cf5488.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
