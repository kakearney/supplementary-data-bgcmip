netcdf CFS-atmos-northPacific-Uwind-2016 {
dimensions:
	wind_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Mon Oct 31 11:55:52 2022: ncks -F -O -d wind_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2016/roms-cfs-atmos-Uwind-2016.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Uwind-2016.nc\n",
			"Mon Sep 10 13:42:58 2018: Time overhang added\n",
			"Mon Sep 10 13:42:50 2018: ncrcat /tmp/tp14d1e34d_b42d_4608_b484_0994faebbb01.nc frc/roms-cfs-atmos-Uwind-2016.nc /tmp/tp994b6b8d_04fb_4504_a302_f22383d2a430.nc /tmp/tpe0ff667b_3374_4228_8222_1a64d4f06c92.nc\n",
			"Mon Sep 10 13:42:50 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2016.nc /tmp/tp14d1e34d_b42d_4608_b484_0994faebbb01.nc\n",
			"Thu Sep  6 14:16:59 2018: ncks -O -F -d wind_time,2,1449 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2016_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2016.nc\n",
			"04-Oct-2017 18:34:55: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
