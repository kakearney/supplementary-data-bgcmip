netcdf CFS-atmos-northPacific-lwrad-2002 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:34 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2002/roms-cfs-atmos-lwrad-2002.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2002/CFS-atmos-northPacific-lwrad-2002.nc\n",
			"Mon Sep 10 13:47:11 2018: Time overhang added\n",
			"Mon Sep 10 13:47:07 2018: ncrcat /tmp/tpaa5df82f_40b8_44f3_9f87_8dd0d01d351d.nc frc/roms-cfs-atmos-lwrad-2002.nc /tmp/tpa6c44327_0361_4eb0_9187_bf4f488ba023.nc /tmp/tp5c5899b6_1ec9_4d0a_a049_375c76b563d8.nc\n",
			"Mon Sep 10 13:47:07 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2002.nc /tmp/tpaa5df82f_40b8_44f3_9f87_8dd0d01d351d.nc\n",
			"Thu Sep  6 10:54:49 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2002_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2002.nc\n",
			"04-Oct-2017 17:55:34: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
