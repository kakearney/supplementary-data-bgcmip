netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-1992 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 14:33:06 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 14:31:26 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1992/CFS-ocean-Bering10K-N30-bryocn-1992.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1992/CFS-ocean-ESPER-Bering10K-N30-brycarbon-1992.nc\n",
			"Wed Dec 14 01:50:48 2022: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad73.nc <>/final/1992/CFS-ocean-Bering10K-N30-bryocn-1992.nc\n",
			"Wed Dec 14 01:49:45 2022: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad01.nc\n",
			"Wed Dec 14 01:49:45 2022: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1992010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1992pentad01.nc\n",
			"Tue Dec 13 06:23:17 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
