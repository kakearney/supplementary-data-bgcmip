netcdf ini_hindcast_unnested_Bering10K_BIO_BANAS {
dimensions:
	xi_rho = 182 ;
	xi_u = 181 ;
	xi_v = 182 ;
	eta_rho = 258 ;
	eta_u = 258 ;
	eta_v = 257 ;
	s_rho = 30 ;
	ocean_time = UNLIMITED ; // (1 currently)
	s_w = 31 ;
variables:
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 1900-01-01 00:00:00" ;
		ocean_time:calendar = "standard" ;
	double zeta(ocean_time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:unit = "meter" ;
		zeta:time = "ocean_time" ;
		zeta:_FillValue = 1.e+36 ;
	double ubar(ocean_time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:unit = "meter second-1" ;
		ubar:time = "ocean_time" ;
		ubar:_FillValue = 1.e+36 ;
	double vbar(ocean_time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:unit = "meter second-1" ;
		vbar:time = "ocean_time" ;
		vbar:_FillValue = 1.e+36 ;
	double u(ocean_time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:unit = "meter second-1" ;
		u:time = "ocean_time" ;
		u:_FillValue = 1.e+36 ;
	double v(ocean_time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:unit = "meter second-1" ;
		v:time = "ocean_time" ;
		v:_FillValue = 1.e+36 ;
	double temp(ocean_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:unit = "Celsius" ;
		temp:time = "ocean_time" ;
		temp:_FillValue = 1.e+36 ;
	double salt(ocean_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:time = "ocean_time" ;
		salt:_FillValue = 1.e+36 ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching function at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching function at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:unit = "meter" ;
	int Vstretching ;
		Vstretching:long_name = "vertical terrain-following stretching function" ;
	int Vtransform ;
		Vtransform:long_name = "vertical terrain-following transformation equation" ;
	double ageice(ocean_time, eta_rho, xi_rho) ;
		ageice:long_name = "age of the ice" ;
		ageice:unit = "sec" ;
		ageice:time = "ocean_time" ;
		ageice:_FillValue = 1.e+36 ;
	double aice(ocean_time, eta_rho, xi_rho) ;
		aice:long_name = "fraction of cell covered by ice" ;
		aice:time = "ocean_time" ;
		aice:_FillValue = 1.e+36 ;
	double h(ocean_time, eta_rho, xi_rho) ;
		h:long_name = "bathymetry at RHO-points" ;
		h:unit = "meter" ;
		h:time = "ocean_time" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:unit = "meter" ;
	double hice(ocean_time, eta_rho, xi_rho) ;
		hice:long_name = "average ice thickness in cell" ;
		hice:unit = "meter" ;
		hice:time = "ocean_time" ;
		hice:_FillValue = 1.e+36 ;
	double lat_rho(ocean_time, eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:unit = "degree_north" ;
		lat_rho:time = "ocean_time" ;
		lat_rho:standard_name = "latitude" ;
	double lat_u(ocean_time, eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:unit = "degree_north" ;
		lat_u:time = "ocean_time" ;
		lat_u:standard_name = "latitude" ;
	double lat_v(ocean_time, eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:unit = "degree_north" ;
		lat_v:time = "ocean_time" ;
		lat_v:standard_name = "latitude" ;
	double lon_rho(ocean_time, eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:unit = "degree_east" ;
		lon_rho:time = "ocean_time" ;
		lon_rho:standard_name = "longitude" ;
	double lon_u(ocean_time, eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:unit = "degree_east" ;
		lon_u:time = "ocean_time" ;
		lon_u:standard_name = "longitude" ;
	double lon_v(ocean_time, eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:unit = "degree_east" ;
		lon_v:time = "ocean_time" ;
		lon_v:standard_name = "longitude" ;
	double s0mk(ocean_time, eta_rho, xi_rho) ;
		s0mk:long_name = "salinity of molecular sub-layer under ice" ;
		s0mk:time = "ocean_time" ;
		s0mk:_FillValue = 1.e+36 ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
		s_rho:positive = "up" ;
		s_rho:standard_name = "ocean_s_coordinate_g1" ;
		s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
		s_w:positive = "up" ;
		s_w:standard_name = "ocean_s_coordinate_g1" ;
		s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
	double sig11(ocean_time, eta_rho, xi_rho) ;
		sig11:long_name = "internal ice stress 11 component" ;
		sig11:unit = "Newton meter-1" ;
		sig11:time = "ocean_time" ;
		sig11:_FillValue = 1.e+36 ;
	double sig12(ocean_time, eta_rho, xi_rho) ;
		sig12:long_name = "internal ice stress 12 component" ;
		sig12:unit = "Newton meter-1" ;
		sig12:time = "ocean_time" ;
		sig12:_FillValue = 1.e+36 ;
	double sig22(ocean_time, eta_rho, xi_rho) ;
		sig22:long_name = "internal ice stress 22 component" ;
		sig22:unit = "Newton meter-1" ;
		sig22:time = "ocean_time" ;
		sig22:_FillValue = 1.e+36 ;
	double snow_thick(ocean_time, eta_rho, xi_rho) ;
		snow_thick:long_name = "thickness of snow cover" ;
		snow_thick:unit = "meter" ;
		snow_thick:time = "ocean_time" ;
		snow_thick:_FillValue = 1.e+36 ;
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = 0., 1. ;
		spherical:flag_meanings = "0 = Cartesian, 1 = spherical" ;
	double t0mk(ocean_time, eta_rho, xi_rho) ;
		t0mk:long_name = "temperature of molecular sub-layer under ice" ;
		t0mk:unit = "Celsius" ;
		t0mk:time = "ocean_time" ;
		t0mk:_FillValue = 1.e+36 ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	double ti(ocean_time, eta_rho, xi_rho) ;
		ti:long_name = "interior ice temperature" ;
		ti:unit = "Celsius" ;
		ti:time = "ocean_time" ;
		ti:_FillValue = 1.e+36 ;
	double tisrf(ocean_time, eta_rho, xi_rho) ;
		tisrf:long_name = "temperature of ice surface" ;
		tisrf:unit = "Celsius" ;
		tisrf:time = "ocean_time" ;
		tisrf:_FillValue = 1.e+36 ;
	double uice(ocean_time, eta_u, xi_u) ;
		uice:long_name = "u-component of ice velocity" ;
		uice:unit = "meter second-1" ;
		uice:time = "ocean_time" ;
		uice:_FillValue = 1.e+36 ;
	double vice(ocean_time, eta_v, xi_v) ;
		vice:long_name = "v-component of ice velocity" ;
		vice:unit = "meter second-1" ;
		vice:time = "ocean_time" ;
		vice:_FillValue = 1.e+36 ;
	double NH4(ocean_time, s_rho, eta_rho, xi_rho) ;
		NH4:long_name = "ammonium" ;
		NH4:unit = "mmol N m^-3" ;
		NH4:time = "ocean_time" ;
		NH4:_FillValue = 1.e+36 ;
	double NO3(ocean_time, s_rho, eta_rho, xi_rho) ;
		NO3:long_name = "nitrate" ;
		NO3:unit = "mmol N m^-3" ;
		NO3:time = "ocean_time" ;
		NO3:_FillValue = 1.e+36 ;
	double det_large(ocean_time, s_rho, eta_rho, xi_rho) ;
		det_large:long_name = "large detritus (aggregates)" ;
		det_large:unit = "mmol N m^-3" ;
		det_large:time = "ocean_time" ;
		det_large:_FillValue = 1.e+36 ;
	double det_small(ocean_time, s_rho, eta_rho, xi_rho) ;
		det_small:long_name = "small detritus" ;
		det_small:unit = "mmol N m^-3" ;
		det_small:time = "ocean_time" ;
		det_small:_FillValue = 1.e+36 ;
	double microzoo(ocean_time, s_rho, eta_rho, xi_rho) ;
		microzoo:long_name = "microzooplankton" ;
		microzoo:unit = "mmol N m^-3" ;
		microzoo:time = "ocean_time" ;
		microzoo:_FillValue = 1.e+36 ;
	double phyto(ocean_time, s_rho, eta_rho, xi_rho) ;
		phyto:long_name = "phytoplankton" ;
		phyto:unit = "mmol N m^-3" ;
		phyto:time = "ocean_time" ;
		phyto:_FillValue = 1.e+36 ;

// global attributes:
		:type = "INITIALIZATION file" ;
		:history = "Wed Jan 25 11:28:26 2023: ncks -A /gscratch/bumblereem/ROMS_Datasets/initial/INIbgc_BIO_BANAS_Bering10K.nc /gscratch/bumblereem/ROMS_Datasets/initial/ini_hindcast_unnested_Bering10K_BIO_BANAS.nc\n",
			"Wed Jan 25 11:27:21 2023: BGC data added: NO3, PO4, Alk, TIC, O2, SiO4: GLODAPv2.2016b Mapped Climatologies; Fe: Huang et al., 2022 climatology + GOANPZ analytical; Hfree, CO3: GLODAPv2 + CO2sys; producers/consumers: seed value; others: 0\n",
			"Wed Jan 25 11:27:20 2023: File schema created via ini_schema.m" ;
		:history_of_appended_files = "Wed Jan 25 11:28:26 2023: Appended file /gscratch/bumblereem/ROMS_Datasets/initial/INIbgc_BIO_BANAS_Bering10K.nc had following \"history\" attribute:\n",
			"Wed Jan 25 11:27:21 2023: BGC data added: NO3, PO4, Alk, TIC, O2, SiO4: GLODAPv2.2016b Mapped Climatologies; Fe: Huang et al., 2022 climatology + GOANPZ analytical; Hfree, CO3: GLODAPv2 + CO2sys; producers/consumers: seed value; others: 0\n",
			"Wed Jan 25 11:27:20 2023: File schema created via ini_schema.m\n",
			"Wed Jan 25 11:28:25 2023: Appended file /gscratch/bumblereem/ROMS_Datasets/initial/INIice_Bering10K.nc had following \"history\" attribute:\n",
			"Wed Jan 25 11:27:04 2023: Ice varible data added: no-ice conditions following ANA_ICE ICE_BASIN example\n",
			"Wed Jan 25 11:27:02 2023: File schema created via ini_schema.m\n",
			"" ;
		:NCO = "4.6.9" ;
}
