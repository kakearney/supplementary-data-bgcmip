netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2015 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 16:33:21 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:30:42 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2015/CFS-ocean-NEP-N30-bryocn-2015.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2015/CFS-ocean-ESPER-NEP-N30-brycarbon-2015.nc\n",
			"Mon Jan  9 23:25:59 2023: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad73.nc <>/final/2015/CFS-ocean-NEP-N30-bryocn-2015.nc\n",
			"Mon Jan  9 23:23:18 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad01.nc\n",
			"Mon Jan  9 23:23:16 2023: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad01.nc\n",
			"Mon Jan  9 23:23:14 2023: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2015010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2015pentad01.nc\n",
			"Mon Jan 09 10:14:31 2023: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
