netcdf INIocean_CFS19900115_NEP {
dimensions:
	xi_rho = 226 ;
	xi_u = 225 ;
	xi_v = 226 ;
	eta_rho = 642 ;
	eta_u = 642 ;
	eta_v = 641 ;
	s_rho = 30 ;
	ocean_time = UNLIMITED ; // (1 currently)
variables:
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 1900-01-01 00:00:00" ;
		ocean_time:calendar = "standard" ;
	double zeta(ocean_time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:unit = "meter" ;
		zeta:time = "ocean_time" ;
		zeta:_FillValue = 1.e+36 ;
	double ubar(ocean_time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:unit = "meter second-1" ;
		ubar:time = "ocean_time" ;
		ubar:_FillValue = 1.e+36 ;
	double vbar(ocean_time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:unit = "meter second-1" ;
		vbar:time = "ocean_time" ;
		vbar:_FillValue = 1.e+36 ;
	double u(ocean_time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:unit = "meter second-1" ;
		u:time = "ocean_time" ;
		u:_FillValue = 1.e+36 ;
	double v(ocean_time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:unit = "meter second-1" ;
		v:time = "ocean_time" ;
		v:_FillValue = 1.e+36 ;
	double temp(ocean_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:unit = "Celsius" ;
		temp:time = "ocean_time" ;
		temp:_FillValue = 1.e+36 ;
	double salt(ocean_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:time = "ocean_time" ;
		salt:_FillValue = 1.e+36 ;

// global attributes:
		:type = "INITIALIZATION file" ;
		:history = "Wed Jan 25 11:28:02 2023: File schema created via ini_schema.m" ;
}
