netcdf CFS-atmos-northPacific-Tair-2015 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:43:34 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2015/roms-cfs-atmos-Tair-2015.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Tair-2015.nc\n",
			"Mon Sep 10 13:39:45 2018: Time overhang added\n",
			"Mon Sep 10 13:39:38 2018: ncrcat /tmp/tp3d69e1a0_7f3f_44f4_bfa3_915dc2aae36b.nc frc/roms-cfs-atmos-Tair-2015.nc /tmp/tpddcb9fd1_3e90_4a8f_8185_88508d6906f6.nc /tmp/tp35965ead_1fd4_4b6b_bf8d_84b172fbddfe.nc\n",
			"Mon Sep 10 13:39:37 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2015.nc /tmp/tp3d69e1a0_7f3f_44f4_bfa3_915dc2aae36b.nc\n",
			"Thu Sep  6 13:41:11 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2015.nc\n",
			"Thu Sep  6 13:39:12 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2015_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2015.nc\n",
			"04-Oct-2017 18:28:54: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
