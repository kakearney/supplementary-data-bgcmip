netcdf CFS-atmos-northPacific-swrad-2016 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	srf_time = UNLIMITED ; // (364 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Mon Oct 31 12:07:21 2022: ncks -F -O -d srf_time,2,365 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2016/roms-cfs-atmos-swrad-2016.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-swrad-2016.nc\n",
			"Mon Sep 10 14:04:38 2018: Time overhang added\n",
			"Mon Sep 10 14:04:35 2018: ncrcat /tmp/tp26316481_50fc_40c7_b175_2c14846ac493.nc frc/roms-cfs-atmos-swrad-2016.nc /tmp/tp5a774eb5_ed20_403f_be86_87aae997a9c6.nc /tmp/tp2a549242_0517_40f5_a220_1337f8986317.nc\n",
			"Mon Sep 10 14:04:35 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-2016.nc /tmp/tp26316481_50fc_40c7_b175_2c14846ac493.nc\n",
			"Thu Sep  6 14:16:35 2018: ncks -O -F -d srf_time,2,365 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2016_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-2016.nc\n",
			"04-Oct-2017 18:34:47: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
