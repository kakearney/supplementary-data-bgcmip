netcdf CFS-atmos-northPacific-lwrad-1996 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1464 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:42:31 2022: ncks -F -O -d lrf_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1996/roms-cfs-atmos-lwrad-1996.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1996/CFS-atmos-northPacific-lwrad-1996.nc\n",
			"Mon Sep 10 13:46:37 2018: Time overhang added\n",
			"Mon Sep 10 13:46:33 2018: ncrcat /tmp/tp7c47faf0_652a_4255_ba32_8ce93ddda977.nc frc/roms-cfs-atmos-lwrad-1996.nc /tmp/tpc0ce6171_fc54_4bff_ae6a_09e8aa397c4d.nc /tmp/tp055c567d_8040_44a5_8447_dbe1b09d6f30.nc\n",
			"Mon Sep 10 13:46:33 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-1996.nc /tmp/tp7c47faf0_652a_4255_ba32_8ce93ddda977.nc\n",
			"Thu Sep  6 09:59:55 2018: ncks -O -F -d lrf_time,2,1465 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1996_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-1996.nc\n",
			"04-Oct-2017 17:40:19: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
