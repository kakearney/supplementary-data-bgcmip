netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-2009 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:59:38 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 15:57:53 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2009/CFS-ocean-Bering10K-N30-bryocn-2009.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2009/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2009.nc\n",
			"Fri Jan  6 09:20:46 2023: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad73.nc <>/final/2009/CFS-ocean-Bering10K-N30-bryocn-2009.nc\n",
			"Fri Jan  6 09:19:30 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad01.nc\n",
			"Fri Jan  6 09:19:30 2023: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad01.nc\n",
			"Fri Jan  6 09:19:30 2023: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2009010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2009pentad01.nc\n",
			"Thu Jan 05 20:03:49 2023: CFS data added\n",
			"Tue Dec 20 15:09:11 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
