netcdf CFS-atmos-northPacific-Uwind-2012 {
dimensions:
	wind_time = UNLIMITED ; // (1464 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:14:46 2022: ncks -F -O -d wind_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2012/roms-cfs-atmos-Uwind-2012.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Uwind-2012.nc\n",
			"Mon Sep 10 13:42:09 2018: Time overhang added\n",
			"Mon Sep 10 13:42:01 2018: ncrcat /tmp/tpd6fa937c_2463_4cdd_8167_bf651bec0d23.nc frc/roms-cfs-atmos-Uwind-2012.nc /tmp/tp29edc1da_b01b_4bed_97f4_22cddafe0009.nc /tmp/tp17815e28_1201_4d4c_9c7d_960272e76640.nc\n",
			"Mon Sep 10 13:42:01 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2012.nc /tmp/tpd6fa937c_2463_4cdd_8167_bf651bec0d23.nc\n",
			"Thu Sep  6 12:46:43 2018: ncks -O -F -d wind_time,2,1465 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2012_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2012.nc\n",
			"04-Oct-2017 18:19:43: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
