netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-2012 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 16:15:13 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:13:28 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2012/CFS-ocean-Bering10K-N30-bryocn-2012.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2012/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2012.nc\n",
			"Sun Jan  8 06:22:44 2023: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad73.nc <>/final/2012/CFS-ocean-Bering10K-N30-bryocn-2012.nc\n",
			"Sun Jan  8 06:21:39 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad01.nc\n",
			"Sun Jan  8 06:21:39 2023: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad01.nc\n",
			"Sun Jan  8 06:21:38 2023: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2012010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2012pentad01.nc\n",
			"Sat Jan 07 16:52:18 2023: CFS data added\n",
			"Tue Dec 20 15:09:11 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
