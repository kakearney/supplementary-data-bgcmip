netcdf CFS-atmos-northPacific-rain-1986 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double rain(rain_time, lat, lon) ;
		rain:missing_value = -1.e+34 ;
		rain:_FillValue = -1.e+34 ;
		rain:time = "rain_time" ;
		rain:coordinates = "lon lat" ;
		rain:long_name = "rainfall" ;
		rain:history = "From roms-cfs-atmos-rain-1986" ;
	double rain_time(rain_time) ;
		rain_time:units = "day since 1900-01-01 00:00:00" ;
		rain_time:time_origin = "01-JAN-1900 00:00:00" ;
		rain_time:axis = "T" ;
		rain_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:20:02 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-rain-1986.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1986/CFS-atmos-northPacific-rain-1986.nc\n",
			"Wed Nov 20 13:49:24 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:49:18 2019: ncrcat /tmp/tpc7896608_a551_4a64_8a58_1747c8c81d4c.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-rain-1986.nc /tmp/tpe0885bc8_d149_477a_b906_26d0579cf67d.nc /tmp/tp6c87f505_ab53_4a95_a29e_d1286c3d6df6.nc\n",
			"Wed Nov 20 13:49:16 2019: ncks -F -d rain_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-rain-1986.nc /tmp/tpc7896608_a551_4a64_8a58_1747c8c81d4c.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
