netcdf CFS-atmos-northPacific-Uwind-2015 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:44:25 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2015/roms-cfs-atmos-Uwind-2015.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Uwind-2015.nc\n",
			"Mon Sep 10 13:42:46 2018: Time overhang added\n",
			"Mon Sep 10 13:42:38 2018: ncrcat /tmp/tp44d38f60_4e33_4056_929e_5ae8d9fe7e7f.nc frc/roms-cfs-atmos-Uwind-2015.nc /tmp/tpd057d87a_9b21_4aa3_8204_4fe660e6bb11.nc /tmp/tpb49a5f5f_848b_498a_be4c_6c74d8b33c19.nc\n",
			"Mon Sep 10 13:42:37 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2015.nc /tmp/tp44d38f60_4e33_4056_929e_5ae8d9fe7e7f.nc\n",
			"Thu Sep  6 13:53:10 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2015_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2015.nc\n",
			"04-Oct-2017 18:31:04: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
