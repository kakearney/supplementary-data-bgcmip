netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2006 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:47:36 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 15:44:27 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2006/CFS-ocean-NEP-N30-bryocn-2006.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2006/CFS-ocean-ESPER-NEP-N30-brycarbon-2006.nc\n",
			"Tue Dec 27 06:37:10 2022: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad73.nc <>/final/2006/CFS-ocean-NEP-N30-bryocn-2006.nc\n",
			"Tue Dec 27 06:35:02 2022: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad01.nc\n",
			"Tue Dec 27 06:35:01 2022: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad01.nc\n",
			"Tue Dec 27 06:35:00 2022: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2006010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2006pentad01.nc\n",
			"Mon Dec 26 17:10:24 2022: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
