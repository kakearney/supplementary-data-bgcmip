netcdf CFS-atmos-northPacific-Uwind-2006 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:52:37 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2006/roms-cfs-atmos-Uwind-2006.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2006/CFS-atmos-northPacific-Uwind-2006.nc\n",
			"Mon Sep 10 13:41:24 2018: Time overhang added\n",
			"Mon Sep 10 13:41:20 2018: ncrcat /tmp/tp980683b9_a8d1_47c3_938b_5700d2041847.nc frc/roms-cfs-atmos-Uwind-2006.nc /tmp/tp2bbea24f_1ebf_4583_8db0_14b62ac6da64.nc /tmp/tpe99cac1c_6555_4fd7_9cff_21914c85bb4d.nc\n",
			"Mon Sep 10 13:41:20 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2006.nc /tmp/tp980683b9_a8d1_47c3_938b_5700d2041847.nc\n",
			"Thu Sep  6 11:36:31 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2006_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2006.nc\n",
			"04-Oct-2017 18:04:32: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
