netcdf CFS-atmos-northPacific-Tair-1997 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:14 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1997/roms-cfs-atmos-Tair-1997.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1997/CFS-atmos-northPacific-Tair-1997.nc\n",
			"Mon Sep 10 13:37:38 2018: Time overhang added\n",
			"Mon Sep 10 13:37:35 2018: ncrcat /tmp/tpce32b1bf_f00d_457f_94c4_12f5c51a2d92.nc frc/roms-cfs-atmos-Tair-1997.nc /tmp/tp0878b2f5_3b74_4fe6_a2a5_0bee4e1c8741.nc /tmp/tp2f1f9dfa_9154_445a_bd8e_ad7ab4a27bf6.nc\n",
			"Mon Sep 10 13:37:34 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-1997.nc /tmp/tpce32b1bf_f00d_457f_94c4_12f5c51a2d92.nc\n",
			"Thu Sep  6 10:07:58 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1997.nc\n",
			"Thu Sep  6 10:07:03 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1997_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1997.nc\n",
			"04-Oct-2017 17:41:45: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
