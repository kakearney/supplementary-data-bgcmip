netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2018 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 16:47:51 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:45:13 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2018/CFS-ocean-NEP-N30-bryocn-2018.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2018/CFS-ocean-ESPER-NEP-N30-brycarbon-2018.nc\n",
			"Wed Jan 11 19:31:43 2023: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad73.nc <>/final/2018/CFS-ocean-NEP-N30-bryocn-2018.nc\n",
			"Wed Jan 11 19:29:44 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad01.nc\n",
			"Wed Jan 11 19:29:43 2023: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad01.nc\n",
			"Wed Jan 11 19:29:43 2023: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2018010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2018pentad01.nc\n",
			"Wed Jan 11 02:53:16 2023: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
