netcdf CFS-atmos-northPacific-Uwind-2000 {
dimensions:
	wind_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:49:04 2022: ncks -F -O -d wind_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2000/roms-cfs-atmos-Uwind-2000.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2000/CFS-atmos-northPacific-Uwind-2000.nc\n",
			"Mon Sep 10 13:40:51 2018: Time overhang added\n",
			"Mon Sep 10 13:40:48 2018: ncrcat /tmp/tp18db8202_a45b_4ea1_80a4_c81672d3051d.nc frc/roms-cfs-atmos-Uwind-2000.nc /tmp/tp143f3a1e_1ab0_40fe_835d_e30182e2ebda.nc /tmp/tpfef920a9_d25b_43a5_ab9a_8f25e3052284.nc\n",
			"Mon Sep 10 13:40:48 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2000.nc /tmp/tp18db8202_a45b_4ea1_80a4_c81672d3051d.nc\n",
			"Thu Sep  6 10:37:00 2018: ncks -O -F -d wind_time,2,1465 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2000_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2000.nc\n",
			"04-Oct-2017 17:50:33: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
