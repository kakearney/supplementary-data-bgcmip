netcdf CFS-atmos-northPacific-Tair-1999 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:47:34 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1999/roms-cfs-atmos-Tair-1999.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1999/CFS-atmos-northPacific-Tair-1999.nc\n",
			"Mon Sep 10 13:37:50 2018: Time overhang added\n",
			"Mon Sep 10 13:37:46 2018: ncrcat /tmp/tp8749915e_beaf_4eae_a9a2_213d581285bb.nc frc/roms-cfs-atmos-Tair-1999.nc /tmp/tp5dcb76f7_8903_47f4_b4ee_8431d0fd6d3d.nc /tmp/tp39d27c72_3f3e_4637_ab1e_52c3527090cf.nc\n",
			"Mon Sep 10 13:37:46 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-1999.nc /tmp/tp8749915e_beaf_4eae_a9a2_213d581285bb.nc\n",
			"Thu Sep  6 10:23:18 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1999.nc\n",
			"Thu Sep  6 10:22:13 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1999_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-1999.nc\n",
			"04-Oct-2017 17:46:41: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
