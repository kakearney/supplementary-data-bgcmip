netcdf CFS-atmos-northPacific-Vwind-2015 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:45:14 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2015/roms-cfs-atmos-Vwind-2015.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Vwind-2015.nc\n",
			"Mon Sep 10 13:45:51 2018: Time overhang added\n",
			"Mon Sep 10 13:45:43 2018: ncrcat /tmp/tpc9069053_5953_499e_915f_bccbdd017635.nc frc/roms-cfs-atmos-Vwind-2015.nc /tmp/tp5eaba7ef_8ddd_4bde_98ad_4f287521cc95.nc /tmp/tp6c50133e_a9ee_4860_85df_2d12eb7c467c.nc\n",
			"Mon Sep 10 13:45:42 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2015.nc /tmp/tpc9069053_5953_499e_915f_bccbdd017635.nc\n",
			"Thu Sep  6 13:55:08 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2015_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2015.nc\n",
			"04-Oct-2017 18:31:04: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
