netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-1999 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:09:39 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 15:08:02 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1999/CFS-ocean-Bering10K-N30-bryocn-1999.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1999/CFS-ocean-ESPER-Bering10K-N30-brycarbon-1999.nc\n",
			"Tue Dec 20 12:07:51 2022: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad73.nc <>/final/1999/CFS-ocean-Bering10K-N30-bryocn-1999.nc\n",
			"Tue Dec 20 12:07:08 2022: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad01.nc\n",
			"Tue Dec 20 12:07:08 2022: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-1999010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-1999pentad01.nc\n",
			"Mon Dec 19 20:57:05 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
