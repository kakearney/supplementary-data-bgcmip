netcdf CFS-atmos-northPacific-Pair-2019 {
dimensions:
	pair_time = UNLIMITED ; // (1457 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:missing_value = -1.e+34 ;
		Pair:_FillValue = -1.e+34 ;
		Pair:time = "pair_time" ;
		Pair:coordinates = "lon lat" ;
		Pair:long_name = "atmos pressure" ;
		Pair:history = "From roms-cfs-atmos-Pair-2019" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double pair_time(pair_time) ;
		pair_time:units = "day since 1900-01-01 00:00:00" ;
		pair_time:time_origin = "01-JAN-1900 00:00:00" ;
		pair_time:axis = "T" ;
		pair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:36:01 2022: ncks -F -O -d pair_time,2,1458 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Pair-2019.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Pair-2019.nc\n",
			"Fri Mar 27 16:03:14 2020: Time overhang added to both ends\n",
			"Fri Mar 27 16:03:05 2020: ncrcat /tmp/tp69921814_f4f7_4d23_a4eb_5834b01a9c42.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Pair-2019.nc /tmp/tp9aca2bb7_ef61_4faa_a8a0_6b2de6217bf9.nc /tmp/tpd99286a3_8020_4796_a6c4_98761f62b522.nc\n",
			"Fri Mar 27 16:03:03 2020: ncks -F -d pair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2019/roms-cfs-atmos-Pair-2019.nc /tmp/tp69921814_f4f7_4d23_a4eb_5834b01a9c42.nc\n",
			"FERRET V7.4   4-Mar-20" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
