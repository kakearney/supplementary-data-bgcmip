netcdf CFS-atmos-northPacific-Pair-2006 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:52:17 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2006/roms-cfs-atmos-Pair-2006.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2006/CFS-atmos-northPacific-Pair-2006.nc\n",
			"Mon Sep 10 13:32:39 2018: Time overhang added\n",
			"Mon Sep 10 13:32:35 2018: ncrcat /tmp/tp87a12a7e_b040_436d_8469_e058a6e72238.nc frc/roms-cfs-atmos-Pair-2006.nc /tmp/tpeea1320b_a3ce_44e5_8c4f_f5e9cf7ae847.nc /tmp/tp52b42f29_183d_46f6_bc20_d26556e91cb1.nc\n",
			"Mon Sep 10 13:32:35 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2006.nc /tmp/tp87a12a7e_b040_436d_8469_e058a6e72238.nc\n",
			"Thu Sep  6 11:29:45 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2006.nc\n",
			"Thu Sep  6 11:28:29 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2006_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2006.nc\n",
			"04-Oct-2017 18:03:25: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
