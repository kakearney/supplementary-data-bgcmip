netcdf CFS-atmos-northPacific-Pair-2011 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:02:21 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2011/roms-cfs-atmos-Pair-2011.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Pair-2011.nc\n",
			"Thu Sep 13 10:47:33 2018: Time overhang added\n",
			"Thu Sep 13 10:47:26 2018: ncrcat /tmp/tp89ca3036_bb2d_4046_a62e_b23fdbb72413.nc frc/roms-cfs-atmos-Pair-2011.nc /tmp/tpfc8f6a89_a493_4d40_a7d3_6095e9dcf1cb.nc /tmp/tp151f6dd8_749b_4111_ac66_1f8a18e98dc8.nc\n",
			"Thu Sep 13 10:47:24 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2011.nc /tmp/tp89ca3036_bb2d_4046_a62e_b23fdbb72413.nc\n",
			"Thu Sep 13 10:40:25 2018: ncrename -d air_time,pair_time -v air_time,pair_time ./frc/roms-cfs-atmos-Pair-2011.nc\n",
			"Thu Sep 13 10:40:15 2018: ncks -O -F -d air_time,2,1461 -v Pair ./frc/Old/corecfs_2011_air.nc ./frc/roms-cfs-atmos-Pair-2011.nc\n",
			"04-Oct-2017 18:13:26: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
