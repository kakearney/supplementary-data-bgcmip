netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-1998 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:07:38 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 15:04:39 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1998/CFS-ocean-NEP-N30-bryocn-1998.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/1998/CFS-ocean-ESPER-NEP-N30-brycarbon-1998.nc\n",
			"Mon Dec 19 20:55:59 2022: ncrcat -O <>/final/1998/CFS-ocean-NEP-N30-bryocn-1998.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad73.nc <>/final/1998/CFS-ocean-NEP-N30-bryocn-1998.nc\n",
			"Mon Dec 19 10:58:02 2022: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad58.nc <>/final/1998/CFS-ocean-NEP-N30-bryocn-1998.nc\n",
			"Mon Dec 19 10:57:19 2022: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad01.nc\n",
			"Mon Dec 19 10:57:18 2022: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1998010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1998pentad01.nc\n",
			"Sat Dec 17 02:36:24 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
