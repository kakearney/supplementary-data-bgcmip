netcdf CFS-atmos-northPacific-Tair-1991 {
dimensions:
	tair_time = UNLIMITED ; // (1459 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:missing_value = -1.e+34 ;
		Tair:_FillValue = -1.e+34 ;
		Tair:time = "tair_time" ;
		Tair:coordinates = "lon lat" ;
		Tair:height_above_ground = 2.f ;
		Tair:long_name = "surface air temperature" ;
		Tair:history = "From roms-cfs-atmos-Tair-1991" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double tair_time(tair_time) ;
		tair_time:units = "day since 1900-01-01 00:00:00" ;
		tair_time:time_origin = "01-JAN-1900 00:00:00" ;
		tair_time:axis = "T" ;
		tair_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:26:13 2022: ncks -F -O -d tair_time,2,1460 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Tair-1991.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1991/CFS-atmos-northPacific-Tair-1991.nc\n",
			"Wed Nov 20 13:58:51 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:58:47 2019: ncrcat /tmp/tpd60aa12e_72eb_43fc_a1f1_5db8a860f2b8.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Tair-1991.nc /tmp/tp15f68227_f1bd_489a_b2d5_9b64c6dedb91.nc /tmp/tp856d7f7f_62de_412b_9dc2_9ac90eeeffe5.nc\n",
			"Wed Nov 20 13:58:46 2019: ncks -F -d tair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Tair-1991.nc /tmp/tpd60aa12e_72eb_43fc_a1f1_5db8a860f2b8.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
