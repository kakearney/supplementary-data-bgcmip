netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2000 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:17:27 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 15:14:32 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2000/CFS-ocean-NEP-N30-bryocn-2000.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2000/CFS-ocean-ESPER-NEP-N30-brycarbon-2000.nc\n",
			"Sat Dec 24 00:51:36 2022: ncrcat -O <>/final/2000/CFS-ocean-NEP-N30-bryocn-2000.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad73.nc <>/final/2000/CFS-ocean-NEP-N30-bryocn-2000.nc\n",
			"Wed Dec 21 13:57:09 2022: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad07.nc <>/final/2000/CFS-ocean-NEP-N30-bryocn-2000.nc\n",
			"Wed Dec 21 13:57:05 2022: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad01.nc\n",
			"Wed Dec 21 13:57:04 2022: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2000010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2000pentad01.nc\n",
			"Tue Dec 20 12:08:46 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
