netcdf CFS-atmos-northPacific-Uwind-1997 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:20 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1997/roms-cfs-atmos-Uwind-1997.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1997/CFS-atmos-northPacific-Uwind-1997.nc\n",
			"Mon Sep 10 13:40:35 2018: Time overhang added\n",
			"Mon Sep 10 13:40:31 2018: ncrcat /tmp/tp20d981d2_d53a_45c5_a2c1_5490f9a2e22b.nc frc/roms-cfs-atmos-Uwind-1997.nc /tmp/tp03cd03a4_f6fc_4ae6_ab25_b1550d757bd7.nc /tmp/tp7510d9e8_7af9_42d5_b210_53b7e98acf6a.nc\n",
			"Mon Sep 10 13:40:31 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-1997.nc /tmp/tp20d981d2_d53a_45c5_a2c1_5490f9a2e22b.nc\n",
			"Thu Sep  6 10:11:30 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1997_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-1997.nc\n",
			"04-Oct-2017 17:43:05: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
