netcdf CFS-atmos-northPacific-Tair-2003 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:17:02 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2003/roms-cfs-atmos-Tair-2003.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2003/CFS-atmos-northPacific-Tair-2003.nc\n",
			"Mon Sep 10 13:38:12 2018: Time overhang added\n",
			"Mon Sep 10 13:38:08 2018: ncrcat /tmp/tp2cd13607_fb38_47b5_8679_808622733f25.nc frc/roms-cfs-atmos-Tair-2003.nc /tmp/tp171b8b03_51d6_4fbb_a852_399cf6572b67.nc /tmp/tp5c40dd7b_06cc_4a5d_a3ce_bb76ffa5c3b9.nc\n",
			"Mon Sep 10 13:38:08 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2003.nc /tmp/tp2cd13607_fb38_47b5_8679_808622733f25.nc\n",
			"Thu Sep  6 11:01:49 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2003.nc\n",
			"Thu Sep  6 11:00:36 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2003_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2003.nc\n",
			"04-Oct-2017 17:57:09: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
