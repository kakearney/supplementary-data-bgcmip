netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-2017 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 16:40:08 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:38:34 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2017/CFS-ocean-Bering10K-N30-bryocn-2017.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2017/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2017.nc\n",
			"Wed Jan 11 02:52:24 2023: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad73.nc <>/final/2017/CFS-ocean-Bering10K-N30-bryocn-2017.nc\n",
			"Wed Jan 11 02:51:14 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad01.nc\n",
			"Wed Jan 11 02:51:13 2023: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad01.nc\n",
			"Wed Jan 11 02:51:13 2023: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2017010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2017pentad01.nc\n",
			"Tue Jan 10 12:58:54 2023: CFS data added\n",
			"Tue Dec 20 15:09:11 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
