netcdf CFS-ocean-NEP-N30-bryocn-1993 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	xi_rho = 226 ;
	xi_u = 225 ;
	xi_v = 226 ;
	s_rho = 30 ;
	eta_rho = 642 ;
	eta_u = 642 ;
	eta_v = 641 ;
variables:
	double bry_time(bry_time) ;
		bry_time:standard_name = "time" ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:axis = "T" ;
	double zeta_south(bry_time, xi_rho) ;
		zeta_south:long_name = "free-surface, southern boundary condition" ;
		zeta_south:_FillValue = -999999. ;
		zeta_south:missing_value = -999999. ;
		zeta_south:unit = "meter" ;
		zeta_south:time = "bry_time" ;
		zeta_south:cell_methods = "bry_time: mean" ;
	double ubar_south(bry_time, xi_u) ;
		ubar_south:long_name = "vertically integrated u-momentum component, southern boundary condition" ;
		ubar_south:_FillValue = -999999. ;
		ubar_south:missing_value = -999999. ;
		ubar_south:unit = "meter second-1" ;
		ubar_south:time = "bry_time" ;
		ubar_south:cell_methods = "bry_time: mean" ;
	double vbar_south(bry_time, xi_v) ;
		vbar_south:long_name = "vertically integrated v-momentum component, southern boundary condition" ;
		vbar_south:_FillValue = -999999. ;
		vbar_south:missing_value = -999999. ;
		vbar_south:unit = "meter second-1" ;
		vbar_south:time = "bry_time" ;
		vbar_south:cell_methods = "bry_time: mean" ;
	double u_south(bry_time, s_rho, xi_u) ;
		u_south:long_name = "u-momentum component, southern boundary condition" ;
		u_south:_FillValue = -999999. ;
		u_south:missing_value = -999999. ;
		u_south:unit = "meter second-1" ;
		u_south:time = "bry_time" ;
		u_south:cell_methods = "bry_time: mean" ;
	double v_south(bry_time, s_rho, xi_v) ;
		v_south:long_name = "v-momentum component, southern boundary condition" ;
		v_south:_FillValue = -999999. ;
		v_south:missing_value = -999999. ;
		v_south:unit = "meter second-1" ;
		v_south:time = "bry_time" ;
		v_south:cell_methods = "bry_time: mean" ;
	double temp_south(bry_time, s_rho, xi_rho) ;
		temp_south:long_name = "potential temperature, southern boundary condition" ;
		temp_south:_FillValue = -999999. ;
		temp_south:missing_value = -999999. ;
		temp_south:unit = "Celsius" ;
		temp_south:time = "bry_time" ;
		temp_south:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:_FillValue = -999999. ;
		salt_south:missing_value = -999999. ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double zeta_west(bry_time, eta_rho) ;
		zeta_west:long_name = "free-surface, western boundary condition" ;
		zeta_west:_FillValue = -999999. ;
		zeta_west:missing_value = -999999. ;
		zeta_west:unit = "meter" ;
		zeta_west:time = "bry_time" ;
		zeta_west:cell_methods = "bry_time: mean" ;
	double ubar_west(bry_time, eta_u) ;
		ubar_west:long_name = "vertically integrated u-momentum component, western boundary condition" ;
		ubar_west:_FillValue = -999999. ;
		ubar_west:missing_value = -999999. ;
		ubar_west:unit = "meter second-1" ;
		ubar_west:time = "bry_time" ;
		ubar_west:cell_methods = "bry_time: mean" ;
	double vbar_west(bry_time, eta_v) ;
		vbar_west:long_name = "vertically integrated v-momentum component, western boundary condition" ;
		vbar_west:_FillValue = -999999. ;
		vbar_west:missing_value = -999999. ;
		vbar_west:unit = "meter second-1" ;
		vbar_west:time = "bry_time" ;
		vbar_west:cell_methods = "bry_time: mean" ;
	double u_west(bry_time, s_rho, eta_u) ;
		u_west:long_name = "u-momentum component, western boundary condition" ;
		u_west:_FillValue = -999999. ;
		u_west:missing_value = -999999. ;
		u_west:unit = "meter second-1" ;
		u_west:time = "bry_time" ;
		u_west:cell_methods = "bry_time: mean" ;
	double v_west(bry_time, s_rho, eta_v) ;
		v_west:long_name = "v-momentum component, western boundary condition" ;
		v_west:_FillValue = -999999. ;
		v_west:missing_value = -999999. ;
		v_west:unit = "meter second-1" ;
		v_west:time = "bry_time" ;
		v_west:cell_methods = "bry_time: mean" ;
	double temp_west(bry_time, s_rho, eta_rho) ;
		temp_west:long_name = "potential temperature, western boundary condition" ;
		temp_west:_FillValue = -999999. ;
		temp_west:missing_value = -999999. ;
		temp_west:unit = "Celsius" ;
		temp_west:time = "bry_time" ;
		temp_west:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:_FillValue = -999999. ;
		salt_west:missing_value = -999999. ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double zeta_east(bry_time, eta_rho) ;
		zeta_east:long_name = "free-surface, eastern boundary condition" ;
		zeta_east:_FillValue = -999999. ;
		zeta_east:missing_value = -999999. ;
		zeta_east:unit = "meter" ;
		zeta_east:time = "bry_time" ;
		zeta_east:cell_methods = "bry_time: mean" ;
	double ubar_east(bry_time, eta_u) ;
		ubar_east:long_name = "vertically integrated u-momentum component, eastern boundary condition" ;
		ubar_east:_FillValue = -999999. ;
		ubar_east:missing_value = -999999. ;
		ubar_east:unit = "meter second-1" ;
		ubar_east:time = "bry_time" ;
		ubar_east:cell_methods = "bry_time: mean" ;
	double vbar_east(bry_time, eta_v) ;
		vbar_east:long_name = "vertically integrated v-momentum component, eastern boundary condition" ;
		vbar_east:_FillValue = -999999. ;
		vbar_east:missing_value = -999999. ;
		vbar_east:unit = "meter second-1" ;
		vbar_east:time = "bry_time" ;
		vbar_east:cell_methods = "bry_time: mean" ;
	double u_east(bry_time, s_rho, eta_u) ;
		u_east:long_name = "u-momentum component, eastern boundary condition" ;
		u_east:_FillValue = -999999. ;
		u_east:missing_value = -999999. ;
		u_east:unit = "meter second-1" ;
		u_east:time = "bry_time" ;
		u_east:cell_methods = "bry_time: mean" ;
	double v_east(bry_time, s_rho, eta_v) ;
		v_east:long_name = "v-momentum component, eastern boundary condition" ;
		v_east:_FillValue = -999999. ;
		v_east:missing_value = -999999. ;
		v_east:unit = "meter second-1" ;
		v_east:time = "bry_time" ;
		v_east:cell_methods = "bry_time: mean" ;
	double temp_east(bry_time, s_rho, eta_rho) ;
		temp_east:long_name = "potential temperature, eastern boundary condition" ;
		temp_east:_FillValue = -999999. ;
		temp_east:missing_value = -999999. ;
		temp_east:unit = "Celsius" ;
		temp_east:time = "bry_time" ;
		temp_east:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:_FillValue = -999999. ;
		salt_east:missing_value = -999999. ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.1.0 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:type = "BOUNDARY file" ;
		:history = "Fri Sep 22 16:55:24 2023: cdo setmissval,-999999 CFS/1993/CFS-ocean-NEP-N30-bryocn-1993.nc test.nc\n",
			"Fri Sep 22 16:38:03 2023: cdo setmissval,nan CFS/1993/CFS-ocean-NEP-N30-bryocn-1993.nc test.nc\n",
			"Wed Dec 14 19:32:51 2022: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad73.nc <>/final/1993/CFS-ocean-NEP-N30-bryocn-1993.nc\n",
			"Wed Dec 14 19:31:27 2022: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad01.nc\n",
			"Wed Dec 14 19:31:27 2022: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-1993010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-1993pentad01.nc\n",
			"Wed Dec 14 01:51:50 2022: CFS data added\n",
			"Fri Dec 09 10:05:18 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
		:CDO = "Climate Data Operators version 2.1.0 (https://mpimet.mpg.de/cdo)" ;
}
