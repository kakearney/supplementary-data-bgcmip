netcdf CFS-atmos-northPacific-swrad-2013 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	srf_time = UNLIMITED ; // (364 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:30:39 2022: ncks -F -O -d srf_time,2,365 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2013/roms-cfs-atmos-swrad-2013.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-swrad-2013.nc\n",
			"Mon Sep 10 14:04:25 2018: Time overhang added\n",
			"Mon Sep 10 14:04:23 2018: ncrcat /tmp/tpaaf3d27e_d35a_4d62_a697_23cc09591ab7.nc frc/roms-cfs-atmos-swrad-2013.nc /tmp/tp21841ac1_a250_4cfb_b039_4b9937102130.nc /tmp/tpb4679311_427e_40d0_a392_afa0110602f9.nc\n",
			"Mon Sep 10 14:04:22 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-2013.nc /tmp/tpaaf3d27e_d35a_4d62_a697_23cc09591ab7.nc\n",
			"Thu Sep  6 13:06:44 2018: ncks -O -F -d srf_time,2,365 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2013_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-2013.nc\n",
			"04-Oct-2017 18:23:24: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
