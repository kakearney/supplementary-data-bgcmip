netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2011 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 16:13:05 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:10:02 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2011/CFS-ocean-NEP-N30-bryocn-2011.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2011/CFS-ocean-ESPER-NEP-N30-brycarbon-2011.nc\n",
			"Sat Jan  7 16:50:02 2023: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad73.nc <>/final/2011/CFS-ocean-NEP-N30-bryocn-2011.nc\n",
			"Sat Jan  7 16:47:50 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad01.nc\n",
			"Sat Jan  7 16:47:50 2023: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad01.nc\n",
			"Sat Jan  7 16:47:49 2023: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2011010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2011pentad01.nc\n",
			"Sat Jan 07 03:20:09 2023: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
