netcdf ini_hindcastloop2_BIO_COBALT {
dimensions:
	ocean_time = UNLIMITED ; // (1 currently)
	s_w = 31 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
	tracer = 31 ;
	s_rho = 30 ;
	boundary = 4 ;
	eta_u = 258 ;
	xi_u = 181 ;
	eta_v = 257 ;
	xi_v = 182 ;
variables:
	float AKs(ocean_time, s_w, eta_rho, xi_rho) ;
		AKs:long_name = "salinity vertical diffusion coefficient" ;
		AKs:units = "meter2 second-1" ;
		AKs:time = "ocean_time" ;
		AKs:grid = "grid" ;
		AKs:location = "face" ;
		AKs:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKs:field = "AKs, scalar, series" ;
	float AKt(ocean_time, s_w, eta_rho, xi_rho) ;
		AKt:long_name = "temperature vertical diffusion coefficient" ;
		AKt:units = "meter2 second-1" ;
		AKt:time = "ocean_time" ;
		AKt:grid = "grid" ;
		AKt:location = "face" ;
		AKt:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKt:field = "AKt, scalar, series" ;
	float AKv(ocean_time, s_w, eta_rho, xi_rho) ;
		AKv:long_name = "vertical viscosity coefficient" ;
		AKv:units = "meter2 second-1" ;
		AKv:time = "ocean_time" ;
		AKv:grid = "grid" ;
		AKv:location = "face" ;
		AKv:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKv:field = "AKv, scalar, series" ;
	double Akt_bak(tracer) ;
		Akt_bak:long_name = "background vertical mixing coefficient for tracers" ;
		Akt_bak:units = "meter2 second-1" ;
	double Akv_bak ;
		Akv_bak:long_name = "background vertical mixing coefficient for momentum" ;
		Akv_bak:units = "meter2 second-1" ;
	int BioIter ;
		BioIter:long_name = "number of iterations to achieve convergence" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
		Cs_r:field = "Cs_r, scalar" ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
		Cs_w:field = "Cs_w, scalar" ;
	double FSobc_in(boundary) ;
		FSobc_in:long_name = "free-surface inflow, nudging inverse time scale" ;
		FSobc_in:units = "second-1" ;
	double FSobc_out(boundary) ;
		FSobc_out:long_name = "free-surface outflow, nudging inverse time scale" ;
		FSobc_out:units = "second-1" ;
	double Falpha ;
		Falpha:long_name = "Power-law shape barotropic filter parameter" ;
	double Fbeta ;
		Fbeta:long_name = "Power-law shape barotropic filter parameter" ;
	double Fgamma ;
		Fgamma:long_name = "Power-law shape barotropic filter parameter" ;
	float Hsbl(ocean_time, eta_rho, xi_rho) ;
		Hsbl:long_name = "depth of oceanic surface boundary layer" ;
		Hsbl:units = "meter" ;
		Hsbl:time = "ocean_time" ;
		Hsbl:grid = "grid" ;
		Hsbl:location = "face" ;
		Hsbl:coordinates = "lon_rho lat_rho ocean_time" ;
		Hsbl:field = "Hsbl, scalar, series" ;
		Hsbl:_FillValue = 1.e+37f ;
	int Lm2CLM ;
		Lm2CLM:long_name = "2D momentum climatology processing switch" ;
		Lm2CLM:flag_values = 0, 1 ;
		Lm2CLM:flag_meanings = ".FALSE. .TRUE." ;
	int Lm3CLM ;
		Lm3CLM:long_name = "3D momentum climatology processing switch" ;
		Lm3CLM:flag_values = 0, 1 ;
		Lm3CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeM2CLM ;
		LnudgeM2CLM:long_name = "2D momentum climatology nudging activation switch" ;
		LnudgeM2CLM:flag_values = 0, 1 ;
		LnudgeM2CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeM3CLM ;
		LnudgeM3CLM:long_name = "3D momentum climatology nudging activation switch" ;
		LnudgeM3CLM:flag_values = 0, 1 ;
		LnudgeM3CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeTCLM(tracer) ;
		LnudgeTCLM:long_name = "tracer climatology nudging activation switch" ;
		LnudgeTCLM:flag_values = 0, 1 ;
		LnudgeTCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LsshCLM ;
		LsshCLM:long_name = "sea surface height climatology processing switch" ;
		LsshCLM:flag_values = 0, 1 ;
		LsshCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerCLM(tracer) ;
		LtracerCLM:long_name = "tracer climatology processing switch" ;
		LtracerCLM:flag_values = 0, 1 ;
		LtracerCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerSponge(tracer) ;
		LtracerSponge:long_name = "horizontal diffusivity sponge activation switch" ;
		LtracerSponge:flag_values = 0, 1 ;
		LtracerSponge:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerSrc(tracer) ;
		LtracerSrc:long_name = "tracer point sources and sink activation switch" ;
		LtracerSrc:flag_values = 0, 1 ;
		LtracerSrc:flag_meanings = ".FALSE. .TRUE." ;
	int LuvSponge ;
		LuvSponge:long_name = "horizontal viscosity sponge activation switch" ;
		LuvSponge:flag_values = 0, 1 ;
		LuvSponge:flag_meanings = ".FALSE. .TRUE." ;
	int LuvSrc ;
		LuvSrc:long_name = "momentum point sources and sink activation switch" ;
		LuvSrc:flag_values = 0, 1 ;
		LuvSrc:flag_meanings = ".FALSE. .TRUE." ;
	int LwSrc ;
		LwSrc:long_name = "mass point sources and sink activation switch" ;
		LwSrc:flag_values = 0, 1 ;
		LwSrc:flag_meanings = ".FALSE. .TRUE." ;
	double M2nudg ;
		M2nudg:long_name = "2D momentum nudging/relaxation inverse time scale" ;
		M2nudg:units = "day-1" ;
	double M2obc_in(boundary) ;
		M2obc_in:long_name = "2D momentum inflow, nudging inverse time scale" ;
		M2obc_in:units = "second-1" ;
	double M2obc_out(boundary) ;
		M2obc_out:long_name = "2D momentum outflow, nudging inverse time scale" ;
		M2obc_out:units = "second-1" ;
	double M3nudg ;
		M3nudg:long_name = "3D momentum nudging/relaxation inverse time scale" ;
		M3nudg:units = "day-1" ;
	double M3obc_in(boundary) ;
		M3obc_in:long_name = "3D momentum inflow, nudging inverse time scale" ;
		M3obc_in:units = "second-1" ;
	double M3obc_out(boundary) ;
		M3obc_out:long_name = "3D momentum outflow, nudging inverse time scale" ;
		M3obc_out:units = "second-1" ;
	int NKML ;
		NKML:long_name = "NKML ?" ;
	double P_C_max_Di ;
		P_C_max_Di:long_name = "P_C_max_Di: Phytoplankton light limitation/growth rate" ;
	double P_C_max_Lg ;
		P_C_max_Lg:long_name = "P_C_max_Lg: Phytoplankton light limitation/growth rate" ;
	double P_C_max_Sm ;
		P_C_max_Sm:long_name = "P_C_max_Sm: Phytoplankton light limitation/growth rate" ;
	double RHO_0 ;
		RHO_0:long_name = "sea water density" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double Tnudg(tracer) ;
		Tnudg:long_name = "Tracers nudging/relaxation inverse time scale" ;
		Tnudg:units = "day-1" ;
	double Tnudg_SSS ;
		Tnudg_SSS:long_name = "SSS nudging/relaxation inverse time scale" ;
		Tnudg_SSS:units = "day-1" ;
	double Tobc_in(boundary, tracer) ;
		Tobc_in:long_name = "tracers inflow, nudging inverse time scale" ;
		Tobc_in:units = "second-1" ;
	double Tobc_out(boundary, tracer) ;
		Tobc_out:long_name = "tracers outflow, nudging inverse time scale" ;
		Tobc_out:units = "second-1" ;
	int Vstretching ;
		Vstretching:long_name = "vertical terrain-following stretching function" ;
	int Vtransform ;
		Vtransform:long_name = "vertical terrain-following transformation equation" ;
	double Znudg ;
		Znudg:long_name = "free-surface nudging/relaxation inverse time scale" ;
		Znudg:units = "day-1" ;
	double Zob ;
		Zob:long_name = "bottom roughness" ;
		Zob:units = "meter" ;
	double Zos ;
		Zos:long_name = "surface roughness" ;
		Zos:units = "meter" ;
	double a1_co2 ;
		a1_co2:long_name = "a1_co2 : Compute the Schmidt number of CO2 in seawater" ;
	double a1_o2 ;
		a1_o2:long_name = "a1_o2 : Compute the Schmidt number of O2 in seawater" ;
	double a2_co2 ;
		a2_co2:long_name = "a2_co2 : Compute the Schmidt number of CO2 in seawater" ;
	double a2_o2 ;
		a2_o2:long_name = "a2_o2 : Compute the Schmidt number of O2 in seawater" ;
	double a3_co2 ;
		a3_co2:long_name = "a3_co2 : Compute the Schmidt number of CO2 in seawater" ;
	double a3_o2 ;
		a3_o2:long_name = "a3_o2 : Compute the Schmidt number of O2 in seawater" ;
	double a4_co2 ;
		a4_co2:long_name = "a4_co2 : Compute the Schmidt number of CO2 in seawater" ;
	double a4_o2 ;
		a4_o2:long_name = "a4_o2 : Compute the Schmidt number of O2 in seawater" ;
	double a_0 ;
		a_0:long_name = "a_0 : coefficients for O2 saturation" ;
	double a_1 ;
		a_1:long_name = "a_1 : coefficients for O2 saturation" ;
	double a_2 ;
		a_2:long_name = "a_2 : coefficients for O2 saturation" ;
	double a_3 ;
		a_3:long_name = "a_3 : coefficients for O2 saturation" ;
	double a_4 ;
		a_4:long_name = "a_4 : coefficients for O2 saturation" ;
	double a_5 ;
		a_5:long_name = "a_5 : coefficients for O2 saturation" ;
	float ageice(ocean_time, eta_rho, xi_rho) ;
		ageice:long_name = "age of the ice" ;
		ageice:units = "sec" ;
		ageice:time = "ocean_time" ;
		ageice:grid = "grid" ;
		ageice:location = "face" ;
		ageice:coordinates = "lon_rho lat_rho ocean_time" ;
		ageice:field = "ice age, scalar, series" ;
		ageice:_FillValue = 1.e+37f ;
	double agg_Di ;
		agg_Di:long_name = "agg_Di: Phytoplankton aggregation" ;
	double agg_Lg ;
		agg_Lg:long_name = "agg_Lg: Phytoplankton aggregation" ;
	double agg_Sm ;
		agg_Sm:long_name = "agg_Sm: Phytoplankton aggregation" ;
	float aice(ocean_time, eta_rho, xi_rho) ;
		aice:long_name = "fraction of cell covered by ice" ;
		aice:time = "ocean_time" ;
		aice:grid = "grid" ;
		aice:location = "face" ;
		aice:coordinates = "lon_rho lat_rho ocean_time" ;
		aice:field = "ice concentration, scalar, series" ;
		aice:_FillValue = 1.e+37f ;
	float alk(ocean_time, s_rho, eta_rho, xi_rho) ;
		alk:long_name = "Alkalinity" ;
		alk:units = "mol/kg" ;
		alk:time = "ocean_time" ;
		alk:grid = "grid" ;
		alk:location = "face" ;
		alk:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		alk:field = "alk, scalar, series" ;
		alk:_FillValue = 1.e+37f ;
	double alk_2_n_denit ;
		alk_2_n_denit:long_name = "alk_2_n_denit: Other stoichiometry" ;
	double alpha_Di ;
		alpha_Di:long_name = "alpha_Di: Phytoplankton light limitation/growth rate" ;
	double alpha_Lg ;
		alpha_Lg:long_name = "alpha_Lg: Phytoplankton light limitation/growth rate" ;
	double alpha_Sm ;
		alpha_Sm:long_name = "alpha_Sm: Phytoplankton light limitation/growth rate" ;
	double alpha_fescav ;
		alpha_fescav:long_name = "alpha_fescav: Iron chemistry" ;
	double b_0 ;
		b_0:long_name = "b_0 : coefficients for O2 saturation" ;
	double b_1 ;
		b_1:long_name = "b_1 : coefficients for O2 saturation" ;
	double b_2 ;
		b_2:long_name = "b_2 : coefficients for O2 saturation" ;
	double b_3 ;
		b_3:long_name = "b_3 : coefficients for O2 saturation" ;
	double beta_fescav ;
		beta_fescav:long_name = "beta_fescav: Iron chemistry" ;
	double bresp_Di ;
		bresp_Di:long_name = "bresp_Di: Phytoplankton light limitation/growth rate" ;
	double bresp_Lg ;
		bresp_Lg:long_name = "bresp_Lg: Phytoplankton light limitation/growth rate" ;
	double bresp_Sm ;
		bresp_Sm:long_name = "bresp_Sm: Phytoplankton light limitation/growth rate" ;
	double bresp_bact ;
		bresp_bact:long_name = "bresp_bact: Bacterial bioenergetics" ;
	double bresp_lgz ;
		bresp_lgz:long_name = "bresp_lgz: Zooplankton bioenergetics" ;
	double bresp_mdz ;
		bresp_mdz:long_name = "bresp_mdz: Zooplankton bioenergetics" ;
	double bresp_smz ;
		bresp_smz:long_name = "bresp_smz: Zooplankton bioenergetics" ;
	double c_0 ;
		c_0:long_name = "c_0 : coefficients for O2 saturation" ;
	double c_2_n ;
		c_2_n:long_name = "c_2_n: Other stoichiometry" ;
	double ca_2_n_arag ;
		ca_2_n_arag:long_name = "ca_2_n_arag: Other stoichiometry" ;
	double ca_2_n_calc ;
		ca_2_n_calc:long_name = "ca_2_n_calc: Other stoichiometry" ;
	double caco3_sat_max ;
		caco3_sat_max:long_name = "caco3_sat_max: Other stoichiometry" ;
	float cadet_arag(ocean_time, s_rho, eta_rho, xi_rho) ;
		cadet_arag:long_name = "Detrital CaCO3" ;
		cadet_arag:units = "mol/kg" ;
		cadet_arag:time = "ocean_time" ;
		cadet_arag:grid = "grid" ;
		cadet_arag:location = "face" ;
		cadet_arag:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		cadet_arag:field = "cadet_arag, scalar, series" ;
		cadet_arag:_FillValue = 1.e+37f ;
	float cadet_calc(ocean_time, s_rho, eta_rho, xi_rho) ;
		cadet_calc:long_name = "Detrital CaCO3" ;
		cadet_calc:units = "mol/kg" ;
		cadet_calc:time = "ocean_time" ;
		cadet_calc:grid = "grid" ;
		cadet_calc:location = "face" ;
		cadet_calc:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		cadet_calc:field = "cadet_calc, scalar, series" ;
		cadet_calc:_FillValue = 1.e+37f ;
	float chl(ocean_time, s_rho, eta_rho, xi_rho) ;
		chl:long_name = "Chlorophyll" ;
		chl:units = "ug kg-1" ;
		chl:time = "ocean_time" ;
		chl:grid = "grid" ;
		chl:location = "face" ;
		chl:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		chl:field = "chl, scalar, series" ;
		chl:_FillValue = 1.e+37f ;
	float chu_iw(ocean_time, eta_rho, xi_rho) ;
		chu_iw:long_name = "ice-water momentum transfer coefficient" ;
		chu_iw:units = "meter second-1" ;
		chu_iw:time = "ocean_time" ;
		chu_iw:grid = "grid" ;
		chu_iw:location = "face" ;
		chu_iw:coordinates = "lon_rho lat_rho ocean_time" ;
		chu_iw:field = "transfer coefficient, scalar, series" ;
		chu_iw:_FillValue = 1.e+37f ;
	float co3_ion(ocean_time, s_rho, eta_rho, xi_rho) ;
		co3_ion:long_name = "Carbonate ion" ;
		co3_ion:units = "mol/kg" ;
		co3_ion:time = "ocean_time" ;
		co3_ion:grid = "grid" ;
		co3_ion:location = "face" ;
		co3_ion:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		co3_ion:field = "co3_ion, scalar, series" ;
		co3_ion:_FillValue = 1.e+37f ;
	double coef_hp ;
		coef_hp:long_name = "coef_hp: Parameters for unresolved higher predators" ;
	float dic(ocean_time, s_rho, eta_rho, xi_rho) ;
		dic:long_name = "Dissolved Inorganic Carbon" ;
		dic:units = "mol/kg" ;
		dic:time = "ocean_time" ;
		dic:grid = "grid" ;
		dic:location = "face" ;
		dic:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		dic:field = "dic, scalar, series" ;
		dic:_FillValue = 1.e+37f ;
	double dstart ;
		dstart:long_name = "time stamp assigned to model initilization" ;
		dstart:units = "days since 1900-01-01 00:00:00" ;
		dstart:calendar = "proleptic_gregorian" ;
	double dt ;
		dt:long_name = "size of long time-steps" ;
		dt:units = "second" ;
	double dtfast ;
		dtfast:long_name = "size of short time-steps" ;
		dtfast:units = "second" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	double exu_Di ;
		exu_Di:long_name = "exu_Di: Phytoplankton losses to exudation" ;
	double exu_Lg ;
		exu_Lg:long_name = "exu_Lg: Phytoplankton losses to exudation" ;
	double exu_Sm ;
		exu_Sm:long_name = "exu_Sm: Phytoplankton losses to exudation" ;
	double fe_2_n_max_Di ;
		fe_2_n_max_Di:long_name = "fe_2_n_max_Di: Nutrient Limitation Parameters (phytoplankton)" ;
	double fe_2_n_max_Lg ;
		fe_2_n_max_Lg:long_name = "fe_2_n_max_Lg: Nutrient Limitation Parameters (phytoplankton)" ;
	double fe_2_n_max_Sm ;
		fe_2_n_max_Sm:long_name = "fe_2_n_max_Sm: Nutrient Limitation Parameters (phytoplankton)" ;
	double fe_2_n_sed ;
		fe_2_n_sed:long_name = "fe_2_n_sed: Iron chemistry" ;
	double fe_2_n_upt_fac ;
		fe_2_n_upt_fac:long_name = "fe_2_n_upt_fac: Nutrient Limitation Parameters (phytoplankton)" ;
	double fe_coast ;
		fe_coast:long_name = "fe_coast: Iron chemistry" ;
	float fed(ocean_time, s_rho, eta_rho, xi_rho) ;
		fed:long_name = "Dissolved Iron" ;
		fed:units = "mol/kg" ;
		fed:time = "ocean_time" ;
		fed:grid = "grid" ;
		fed:location = "face" ;
		fed:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		fed:field = "fed, scalar, series" ;
		fed:_FillValue = 1.e+37f ;
	float fedet(ocean_time, s_rho, eta_rho, xi_rho) ;
		fedet:long_name = "Detrital Iron" ;
		fedet:units = "mol/kg" ;
		fedet:time = "ocean_time" ;
		fedet:grid = "grid" ;
		fedet:location = "face" ;
		fedet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		fedet:field = "fedet, scalar, series" ;
		fedet:_FillValue = 1.e+37f ;
	float fedi(ocean_time, s_rho, eta_rho, xi_rho) ;
		fedi:long_name = "Diazotroph Iron" ;
		fedi:units = "mol/kg" ;
		fedi:time = "ocean_time" ;
		fedi:grid = "grid" ;
		fedi:location = "face" ;
		fedi:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		fedi:field = "fedi, scalar, series" ;
		fedi:_FillValue = 1.e+37f ;
	float felg(ocean_time, s_rho, eta_rho, xi_rho) ;
		felg:long_name = "Large Phytoplankton Iron" ;
		felg:units = "mol/kg" ;
		felg:time = "ocean_time" ;
		felg:grid = "grid" ;
		felg:location = "face" ;
		felg:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		felg:field = "felg, scalar, series" ;
		felg:_FillValue = 1.e+37f ;
	double felig_2_don ;
		felig_2_don:long_name = "felig_2_don: Iron chemistry" ;
	double felig_bkg ;
		felig_bkg:long_name = "felig_bkg: Iron chemistry" ;
	float fesm(ocean_time, s_rho, eta_rho, xi_rho) ;
		fesm:long_name = "Small Phytoplankton Iron" ;
		fesm:units = "mol/kg" ;
		fesm:time = "ocean_time" ;
		fesm:grid = "grid" ;
		fesm:location = "face" ;
		fesm:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		fesm:field = "fesm, scalar, series" ;
		fesm:_FillValue = 1.e+37f ;
	double ffe_sed_max ;
		ffe_sed_max:long_name = "ffe_sed_max: Iron chemistry" ;
	double gamma2 ;
		gamma2:long_name = "slipperiness parameter" ;
	double gamma_cadet_arag ;
		gamma_cadet_arag:long_name = "gamma_cadet_arag: Remineralization" ;
	double gamma_cadet_calc ;
		gamma_cadet_calc:long_name = "gamma_cadet_calc: Remineralization" ;
	double gamma_fescav ;
		gamma_fescav:long_name = "gamma_fescav: Iron chemistry" ;
	double gamma_irr_mem ;
		gamma_irr_mem:long_name = "gamma_irr_mem: Phytoplankton light limitation/growth rate" ;
	double gamma_mu_mem ;
		gamma_mu_mem:long_name = "gamma_mu_mem: Phytoplankton aggregation limit rate" ;
	double gamma_ndet ;
		gamma_ndet:long_name = "gamma_ndet: Remineralization" ;
	double gamma_nitrif ;
		gamma_nitrif:long_name = "gamma_nitrif: Nitrification" ;
	double gamma_sidet ;
		gamma_sidet:long_name = "gamma_sidet: Remineralization" ;
	double gamma_sldon ;
		gamma_sldon:long_name = "gamma_sldon: Dissolved Organic Material" ;
	double gamma_sldop ;
		gamma_sldop:long_name = "gamma_sldop: Dissolved Organic Material" ;
	double gamma_srdon ;
		gamma_srdon:long_name = "gamma_srdon: Dissolved Organic Material" ;
	double gamma_srdop ;
		gamma_srdop:long_name = "gamma_srdop: Dissolved Organic Material" ;
	double gge_max_bact ;
		gge_max_bact:long_name = "gge_max_bact: Bacterial bioenergetics" ;
	double gge_max_lgz ;
		gge_max_lgz:long_name = "gge_max_lgz: Zooplankton bioenergetics" ;
	double gge_max_mdz ;
		gge_max_mdz:long_name = "gge_max_mdz: Zooplankton bioenergetics" ;
	double gge_max_smz ;
		gge_max_smz:long_name = "gge_max_smz: Zooplankton bioenergetics" ;
	int grid ;
		grid:cf_role = "grid_topology" ;
		grid:topology_dimension = 2 ;
		grid:node_dimensions = "xi_psi eta_psi" ;
		grid:face_dimensions = "xi_rho: xi_psi (padding: both) eta_rho: eta_psi (padding: both)" ;
		grid:edge1_dimensions = "xi_u: xi_psi eta_u: eta_psi (padding: both)" ;
		grid:edge2_dimensions = "xi_v: xi_psi (padding: both) eta_v: eta_psi" ;
		grid:node_coordinates = "lon_psi lat_psi" ;
		grid:face_coordinates = "lon_rho lat_rho" ;
		grid:edge1_coordinates = "lon_u lat_u" ;
		grid:edge2_coordinates = "lon_v lat_v" ;
		grid:vertical_dimensions = "s_rho: s_w (padding: none)" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	float hice(ocean_time, eta_rho, xi_rho) ;
		hice:long_name = "average ice thickness in cell" ;
		hice:units = "meter" ;
		hice:time = "ocean_time" ;
		hice:grid = "grid" ;
		hice:location = "face" ;
		hice:coordinates = "lon_rho lat_rho ocean_time" ;
		hice:field = "ice thickness, scalar, series" ;
		hice:_FillValue = 1.e+37f ;
	double hp_ipa_bact ;
		hp_ipa_bact:long_name = "hp_ipa_bact: Parameters for unresolved higher predators" ;
	double hp_ipa_det ;
		hp_ipa_det:long_name = "hp_ipa_det: Parameters for unresolved higher predators" ;
	double hp_ipa_diaz ;
		hp_ipa_diaz:long_name = "hp_ipa_diaz: Parameters for unresolved higher predators" ;
	double hp_ipa_lgp ;
		hp_ipa_lgp:long_name = "hp_ipa_lgp: Parameters for unresolved higher predators" ;
	double hp_ipa_lgz ;
		hp_ipa_lgz:long_name = "hp_ipa_lgz: Parameters for unresolved higher predators" ;
	double hp_ipa_mdz ;
		hp_ipa_mdz:long_name = "hp_ipa_mdz: Parameters for unresolved higher predators" ;
	double hp_ipa_smp ;
		hp_ipa_smp:long_name = "hp_ipa_smp: Parameters for unresolved higher predators" ;
	double hp_ipa_smz ;
		hp_ipa_smz:long_name = "hp_ipa_smz: Parameters for unresolved higher predators" ;
	double hp_phi_det ;
		hp_phi_det:long_name = "hp_phi_det: Parameters for unresolved higher predators" ;
	double hp_phi_ldon ;
		hp_phi_ldon:long_name = "hp_phi_ldon: Parameters for unresolved higher predators" ;
	double hp_phi_ldop ;
		hp_phi_ldop:long_name = "hp_phi_ldop: Parameters for unresolved higher predators" ;
	double hp_phi_nh4 ;
		hp_phi_nh4:long_name = "hp_phi_nh4: Parameters for unresolved higher predators" ;
	double hp_phi_po4 ;
		hp_phi_po4:long_name = "hp_phi_po4: Parameters for unresolved higher predators" ;
	double hp_phi_sldon ;
		hp_phi_sldon:long_name = "hp_phi_sldon: Parameters for unresolved higher predators" ;
	double hp_phi_sldop ;
		hp_phi_sldop:long_name = "hp_phi_sldop: Parameters for unresolved higher predators" ;
	double hp_phi_srdon ;
		hp_phi_srdon:long_name = "hp_phi_srdon: Parameters for unresolved higher predators" ;
	double hp_phi_srdop ;
		hp_phi_srdop:long_name = "hp_phi_srdop: Parameters for unresolved higher predators" ;
	float htotal(ocean_time, s_rho, eta_rho, xi_rho) ;
		htotal:long_name = "H+ ion concentration" ;
		htotal:units = "mol/kg" ;
		htotal:time = "ocean_time" ;
		htotal:grid = "grid" ;
		htotal:location = "face" ;
		htotal:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		htotal:field = "htotal, scalar, series" ;
		htotal:_FillValue = 1.e+37f ;
	double htotal_in ;
		htotal_in:long_name = "htotal_in: ?" ;
	double htotal_scale_hi ;
		htotal_scale_hi:long_name = "htotal_scale_hi ?" ;
	double htotal_scale_lo ;
		htotal_scale_lo:long_name = "htotal_scale_lo ?" ;
		htotal_scale_lo:units = "?" ;
	double imax_hp ;
		imax_hp:long_name = "imax_hp: Parameters for unresolved higher predators" ;
	double imax_lgz ;
		imax_lgz:long_name = "imax_lgz: Zooplankton ingestion parameterization and temperature dependence" ;
	double imax_mdz ;
		imax_mdz:long_name = "imax_mdz: Zooplankton ingestion parameterization and temperature dependence" ;
	double imax_smz ;
		imax_smz:long_name = "imax_smz: Zooplankton ingestion parameterization and temperature dependence" ;
	double io_fescav ;
		io_fescav:long_name = "io_fescav: Iron chemistry" ;
	double irr_inhibit ;
		irr_inhibit:long_name = "irr_inhibit: Nitrification" ;
	float irr_mem(ocean_time, s_rho, eta_rho, xi_rho) ;
		irr_mem:long_name = "Irradiance memory" ;
		irr_mem:units = "Watts/m^2" ;
		irr_mem:time = "ocean_time" ;
		irr_mem:grid = "grid" ;
		irr_mem:location = "face" ;
		irr_mem:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		irr_mem:field = "irr_mem, scalar, series" ;
		irr_mem:_FillValue = 1.e+37f ;
	double k_fe_2_n_Di ;
		k_fe_2_n_Di:long_name = "k_fe_2_n_Di: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_fe_2_n_Lg ;
		k_fe_2_n_Lg:long_name = "k_fe_2_n_Lg: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_fe_2_n_Sm ;
		k_fe_2_n_Sm:long_name = "k_fe_2_n_Sm: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_fed_Di ;
		k_fed_Di:long_name = "k_fed_Di: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_fed_Lg ;
		k_fed_Lg:long_name = "k_fed_Lg: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_fed_Sm ;
		k_fed_Sm:long_name = "k_fed_Sm: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_ldon_bact ;
		k_ldon_bact:long_name = "k_ldon_bact: Bacterial growth and uptake parameters" ;
	double k_lith ;
		k_lith:long_name = "k_lith: Remineralization" ;
	double k_n_inhib_Di ;
		k_n_inhib_Di:long_name = "k_n_inhib_Di: Nitrogen fixation inhibition parameters" ;
	double k_nh4_Di ;
		k_nh4_Di:long_name = "k_nh4_Di: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_nh4_Lg ;
		k_nh4_Lg:long_name = "k_nh4_Lg: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_nh4_Sm ;
		k_nh4_Sm:long_name = "k_nh4_Sm: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_no3_Di ;
		k_no3_Di:long_name = "k_no3_Di: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_no3_Lg ;
		k_no3_Lg:long_name = "k_no3_Lg: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_no3_Sm ;
		k_no3_Sm:long_name = "k_no3_Sm: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_no3_denit ;
		k_no3_denit:long_name = "k_no3_denit: Remineralization" ;
	double k_o2 ;
		k_o2:long_name = "k_o2: Remineralization" ;
	double k_po4_Di ;
		k_po4_Di:long_name = "k_po4_Di: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_po4_Lg ;
		k_po4_Lg:long_name = "k_po4_Lg: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_po4_Sm ;
		k_po4_Sm:long_name = "k_po4_Sm: Nutrient Limitation Parameters (phytoplankton)" ;
	double k_sed1 ;
		k_sed1:long_name = "Depth-based attenuation coefficient, factor" ;
		k_sed1:units = "m^-1" ;
	double k_sed2 ;
		k_sed2:long_name = "Depth-based attenuation coefficient, exponent" ;
		k_sed2:units = "unitless" ;
	double k_sio4_Lg ;
		k_sio4_Lg:long_name = "k_sio4_Lg: Nutrient Limitation Parameters (phytoplankton)" ;
	double kappa_eppley ;
		kappa_eppley:long_name = "kappa_eppley: Phytoplankton light limitation/growth rate" ;
	double kfe_eq_lig_hl ;
		kfe_eq_lig_hl:long_name = "kfe_eq_lig_hl: Iron chemistry" ;
	double kfe_eq_lig_ll ;
		kfe_eq_lig_ll:long_name = "kfe_eq_lig_ll: Iron chemistry" ;
	double ki_fescav ;
		ki_fescav:long_name = "ki_fescav: Iron chemistry" ;
	double ki_hp ;
		ki_hp:long_name = "ki_hp: Parameters for unresolved higher predators" ;
	double ki_lgz ;
		ki_lgz:long_name = "ki_lgz: Zooplankton ingestion parameterization and temperature dependence" ;
	double ki_mdz ;
		ki_mdz:long_name = "ki_mdz: Zooplankton ingestion parameterization and temperature dependence" ;
	double ki_smz ;
		ki_smz:long_name = "ki_smz: Zooplankton ingestion parameterization and temperature dependence" ;
	double ktemp_bact ;
		ktemp_bact:long_name = "ktemp_bact: Bacterial growth and uptake parameters" ;
	double ktemp_hp ;
		ktemp_hp:long_name = "ktemp_hp: Parameters for unresolved higher predators" ;
	double ktemp_lgz ;
		ktemp_lgz:long_name = "ktemp_lgz: Zooplankton ingestion parameterization and temperature dependence" ;
	double ktemp_mdz ;
		ktemp_mdz:long_name = "ktemp_mdz: Zooplankton ingestion parameterization and temperature dependence" ;
	double ktemp_smz ;
		ktemp_smz:long_name = "ktemp_smz: Zooplankton ingestion parameterization and temperature dependence" ;
	double ktemp_vir ;
		ktemp_vir:long_name = "ktemp_vir: Phytoplankton and bacterial losses to viruses" ;
	float ldon(ocean_time, s_rho, eta_rho, xi_rho) ;
		ldon:long_name = "labile DON" ;
		ldon:units = "mol/kg" ;
		ldon:time = "ocean_time" ;
		ldon:grid = "grid" ;
		ldon:location = "face" ;
		ldon:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		ldon:field = "ldon, scalar, series" ;
		ldon:_FillValue = 1.e+37f ;
	double lgz_ipa_bact ;
		lgz_ipa_bact:long_name = "lgz_ipa_bact: Zooplankton switching and prey preference parameters" ;
	double lgz_ipa_det ;
		lgz_ipa_det:long_name = "lgz_ipa_det: Zooplankton switching and prey preference parameters" ;
	double lgz_ipa_diaz ;
		lgz_ipa_diaz:long_name = "lgz_ipa_diaz: Zooplankton switching and prey preference parameters" ;
	double lgz_ipa_lgp ;
		lgz_ipa_lgp:long_name = "lgz_ipa_lgp: Zooplankton switching and prey preference parameters" ;
	double lgz_ipa_lgz ;
		lgz_ipa_lgz:long_name = "lgz_ipa_lgz: Zooplankton switching and prey preference parameters" ;
	double lgz_ipa_mdz ;
		lgz_ipa_mdz:long_name = "lgz_ipa_mdz: Zooplankton switching and prey preference parameters" ;
	double lgz_ipa_smp ;
		lgz_ipa_smp:long_name = "lgz_ipa_smp: Zooplankton switching and prey preference parameters" ;
	double lgz_ipa_smz ;
		lgz_ipa_smz:long_name = "lgz_ipa_smz: Zooplankton switching and prey preference parameters" ;
	float lith(ocean_time, s_rho, eta_rho, xi_rho) ;
		lith:long_name = "Lithogenic Aluminosilicate" ;
		lith:units = "g/kg" ;
		lith:time = "ocean_time" ;
		lith:grid = "grid" ;
		lith:location = "face" ;
		lith:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		lith:field = "lith, scalar, series" ;
		lith:_FillValue = 1.e+37f ;
	float lithdet(ocean_time, s_rho, eta_rho, xi_rho) ;
		lithdet:long_name = "lithdet" ;
		lithdet:units = "g/kg" ;
		lithdet:time = "ocean_time" ;
		lithdet:grid = "grid" ;
		lithdet:location = "face" ;
		lithdet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		lithdet:field = "lithdet, scalar, series" ;
		lithdet:_FillValue = 1.e+37f ;
	double mass_2_n ;
		mass_2_n:long_name = "mass_2_n: Stoichiometry" ;
	double mdz_ipa_bact ;
		mdz_ipa_bact:long_name = "mdz_ipa_bact: Zooplankton switching and prey preference parameters" ;
	double mdz_ipa_det ;
		mdz_ipa_det:long_name = "mdz_ipa_det: Zooplankton switching and prey preference parameters" ;
	double mdz_ipa_diaz ;
		mdz_ipa_diaz:long_name = "mdz_ipa_diaz: Zooplankton switching and prey preference parameters" ;
	double mdz_ipa_lgp ;
		mdz_ipa_lgp:long_name = "mdz_ipa_lgp: Zooplankton switching and prey preference parameters" ;
	double mdz_ipa_lgz ;
		mdz_ipa_lgz:long_name = "mdz_ipa_lgz: Zooplankton switching and prey preference parameters" ;
	double mdz_ipa_mdz ;
		mdz_ipa_mdz:long_name = "mdz_ipa_mdz: Zooplankton switching and prey preference parameters" ;
	double mdz_ipa_smp ;
		mdz_ipa_smp:long_name = "mdz_ipa_smp: Zooplankton switching and prey preference parameters" ;
	double mdz_ipa_smz ;
		mdz_ipa_smz:long_name = "mdz_ipa_smz: Zooplankton switching and prey preference parameters" ;
	double mswitch_hp ;
		mswitch_hp:long_name = "mswitch_hp: Parameters for unresolved higher predators" ;
	double mswitch_lgz ;
		mswitch_lgz:long_name = "mswitch_lgz: Zooplankton switching and prey preference parameters" ;
	double mswitch_mdz ;
		mswitch_mdz:long_name = "mswitch_mdz: Zooplankton switching and prey preference parameters" ;
	double mswitch_smz ;
		mswitch_smz:long_name = "mswitch_smz: Zooplankton switching and prey preference parameters" ;
	double mu_max_bact ;
		mu_max_bact:long_name = "mu_max_bact: Bacterial growth and uptake parameters" ;
	float mu_mem_di(ocean_time, s_rho, eta_rho, xi_rho) ;
		mu_mem_di:long_name = "Aggreg memory diatoms" ;
		mu_mem_di:units = "None" ;
		mu_mem_di:time = "ocean_time" ;
		mu_mem_di:grid = "grid" ;
		mu_mem_di:location = "face" ;
		mu_mem_di:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		mu_mem_di:field = "mu_mem_di, scalar, series" ;
		mu_mem_di:_FillValue = 1.e+37f ;
	float mu_mem_lg(ocean_time, s_rho, eta_rho, xi_rho) ;
		mu_mem_lg:long_name = "Aggreg memory large phyto" ;
		mu_mem_lg:units = "None" ;
		mu_mem_lg:time = "ocean_time" ;
		mu_mem_lg:grid = "grid" ;
		mu_mem_lg:location = "face" ;
		mu_mem_lg:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		mu_mem_lg:field = "mu_mem_lg, scalar, series" ;
		mu_mem_lg:_FillValue = 1.e+37f ;
	float mu_mem_sm(ocean_time, s_rho, eta_rho, xi_rho) ;
		mu_mem_sm:long_name = "Aggreg memory small phyto" ;
		mu_mem_sm:units = "None" ;
		mu_mem_sm:time = "ocean_time" ;
		mu_mem_sm:grid = "grid" ;
		mu_mem_sm:location = "face" ;
		mu_mem_sm:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		mu_mem_sm:field = "mu_mem_sm, scalar, series" ;
		mu_mem_sm:_FillValue = 1.e+37f ;
	int nAVG ;
		nAVG:long_name = "number of time-steps between time-averaged records" ;
	int nDIA ;
		nDIA:long_name = "number of time-steps between diagnostic records" ;
	int nHIS ;
		nHIS:long_name = "number of time-steps between history records" ;
	int nRST ;
		nRST:long_name = "number of time-steps between restart records" ;
		nRST:cycle = "only latest two records are maintained" ;
	int nSTA ;
		nSTA:long_name = "number of time-steps between stations records" ;
	double n_2_n_denit ;
		n_2_n_denit:long_name = "n_2_n_denit: Stoichiometry" ;
	float nbact(ocean_time, s_rho, eta_rho, xi_rho) ;
		nbact:long_name = "bacterial" ;
		nbact:units = "mol/kg" ;
		nbact:time = "ocean_time" ;
		nbact:grid = "grid" ;
		nbact:location = "face" ;
		nbact:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		nbact:field = "nbact, scalar, series" ;
		nbact:_FillValue = 1.e+37f ;
	int ndefAVG ;
		ndefAVG:long_name = "number of time-steps between the creation of average files" ;
	int ndefDIA ;
		ndefDIA:long_name = "number of time-steps between the creation of diagnostic files" ;
	int ndefHIS ;
		ndefHIS:long_name = "number of time-steps between the creation of history files" ;
	float ndet(ocean_time, s_rho, eta_rho, xi_rho) ;
		ndet:long_name = "ndet" ;
		ndet:units = "mol/kg" ;
		ndet:time = "ocean_time" ;
		ndet:grid = "grid" ;
		ndet:location = "face" ;
		ndet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		ndet:field = "ndet, scalar, series" ;
		ndet:_FillValue = 1.e+37f ;
	float ndi(ocean_time, s_rho, eta_rho, xi_rho) ;
		ndi:long_name = "Diazotroph Nitrogen" ;
		ndi:units = "mol/kg" ;
		ndi:time = "ocean_time" ;
		ndi:grid = "grid" ;
		ndi:location = "face" ;
		ndi:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		ndi:field = "ndi, scalar, series" ;
		ndi:_FillValue = 1.e+37f ;
	int ndtfast ;
		ndtfast:long_name = "number of short time-steps" ;
	float nh4(ocean_time, s_rho, eta_rho, xi_rho) ;
		nh4:long_name = "Ammonia" ;
		nh4:units = "mol/kg" ;
		nh4:time = "ocean_time" ;
		nh4:grid = "grid" ;
		nh4:location = "face" ;
		nh4:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		nh4:field = "nh4, scalar, series" ;
		nh4:_FillValue = 1.e+37f ;
	double nl_tnu2(tracer) ;
		nl_tnu2:long_name = "nonlinear model Laplacian mixing coefficient for tracers" ;
		nl_tnu2:units = "meter2 second-1" ;
	double nl_visc2 ;
		nl_visc2:long_name = "nonlinear model Laplacian mixing coefficient for momentum" ;
		nl_visc2:units = "meter2 second-1" ;
	float nlg(ocean_time, s_rho, eta_rho, xi_rho) ;
		nlg:long_name = "Large Phytoplankton Nitrogen" ;
		nlg:units = "mol/kg" ;
		nlg:time = "ocean_time" ;
		nlg:grid = "grid" ;
		nlg:location = "face" ;
		nlg:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		nlg:field = "nlg, scalar, series" ;
		nlg:_FillValue = 1.e+37f ;
	float nlgz(ocean_time, s_rho, eta_rho, xi_rho) ;
		nlgz:long_name = "large Zooplankton Nitrogen" ;
		nlgz:units = "mol/kg" ;
		nlgz:time = "ocean_time" ;
		nlgz:grid = "grid" ;
		nlgz:location = "face" ;
		nlgz:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		nlgz:field = "nlgz, scalar, series" ;
		nlgz:_FillValue = 1.e+37f ;
	float nmdz(ocean_time, s_rho, eta_rho, xi_rho) ;
		nmdz:long_name = "Medium-sized zooplankton Nitrogen" ;
		nmdz:units = "mol/kg" ;
		nmdz:time = "ocean_time" ;
		nmdz:grid = "grid" ;
		nmdz:location = "face" ;
		nmdz:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		nmdz:field = "nmdz, scalar, series" ;
		nmdz:_FillValue = 1.e+37f ;
	float no3(ocean_time, s_rho, eta_rho, xi_rho) ;
		no3:long_name = "Nitrate" ;
		no3:units = "mol/kg" ;
		no3:time = "ocean_time" ;
		no3:grid = "grid" ;
		no3:location = "face" ;
		no3:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		no3:field = "no3, scalar, series" ;
		no3:_FillValue = 1.e+37f ;
	float nsm(ocean_time, s_rho, eta_rho, xi_rho) ;
		nsm:long_name = "Small Phytoplankton Nitrogen" ;
		nsm:units = "mol/kg" ;
		nsm:time = "ocean_time" ;
		nsm:grid = "grid" ;
		nsm:location = "face" ;
		nsm:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		nsm:field = "nsm, scalar, series" ;
		nsm:_FillValue = 1.e+37f ;
	float nsmz(ocean_time, s_rho, eta_rho, xi_rho) ;
		nsmz:long_name = "Small Zooplankton Nitrogen" ;
		nsmz:units = "mol/kg" ;
		nsmz:time = "ocean_time" ;
		nsmz:grid = "grid" ;
		nsmz:location = "face" ;
		nsmz:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		nsmz:field = "nsmz, scalar, series" ;
		nsmz:_FillValue = 1.e+37f ;
	double nswitch_hp ;
		nswitch_hp:long_name = "nswitch_hp: Parameters for unresolved higher predators" ;
	double nswitch_lgz ;
		nswitch_lgz:long_name = "nswitch_lgz: Zooplankton switching and prey preference parameters" ;
	double nswitch_mdz ;
		nswitch_mdz:long_name = "nswitch_mdz: Zooplankton switching and prey preference parameters" ;
	double nswitch_smz ;
		nswitch_smz:long_name = "nswitch_smz: Zooplankton switching and prey preference parameters" ;
	int ntimes ;
		ntimes:long_name = "number of long time-steps" ;
	int ntsAVG ;
		ntsAVG:long_name = "starting time-step for accumulation of time-averaged fields" ;
	int ntsDIA ;
		ntsDIA:long_name = "starting time-step for accumulation of diagnostic fields" ;
	float o2(ocean_time, s_rho, eta_rho, xi_rho) ;
		o2:long_name = "Oxygen" ;
		o2:units = "mol/kg" ;
		o2:time = "ocean_time" ;
		o2:grid = "grid" ;
		o2:location = "face" ;
		o2:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		o2:field = "o2, scalar, series" ;
		o2:_FillValue = 1.e+37f ;
	double o2_2_c ;
		o2_2_c:long_name = "o2_2_c: Stoichiometry" ;
	double o2_2_nfix ;
		o2_2_nfix:long_name = "o2_2_nfix: Stoichiometry" ;
	double o2_2_nh4 ;
		o2_2_nh4:long_name = "o2_2_nh4: Stoichiometry" ;
	double o2_2_nitrif ;
		o2_2_nitrif:long_name = "o2_2_nitrif: Stoichiometry" ;
	double o2_2_no3 ;
		o2_2_no3:long_name = "o2_2_no3: Stoichiometry" ;
	double o2_inhib_Di_pow ;
		o2_inhib_Di_pow:long_name = "o2_inhib_Di_pow: Nitrogen fixation inhibition parameters" ;
	double o2_inhib_Di_sat ;
		o2_inhib_Di_sat:long_name = "o2_inhib_Di_sat: Nitrogen fixation inhibition parameters" ;
	double o2_min ;
		o2_min:long_name = "o2_min: Remineralization" ;
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 1900-01-01 00:00:00" ;
		ocean_time:calendar = "proleptic_gregorian" ;
		ocean_time:field = "time, scalar, series" ;
	int p_2_n_static ;
		p_2_n_static:long_name = "p_2_n_static: Other stoichiometry" ;
	double p_2_n_static_Di ;
		p_2_n_static_Di:long_name = "p_2_n_static_Di: Other stoichiometry" ;
	double p_2_n_static_Lg ;
		p_2_n_static_Lg:long_name = "p_2_n_static_Lg: Other stoichiometry" ;
	double p_2_n_static_Sm ;
		p_2_n_static_Sm:long_name = "p_2_n_static_Sm: Other stoichiometry" ;
	double phi_det_lgz ;
		phi_det_lgz:long_name = "phi_det_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_det_mdz ;
		phi_det_mdz:long_name = "phi_det_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_det_smz ;
		phi_det_smz:long_name = "phi_det_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_ldon_lgz ;
		phi_ldon_lgz:long_name = "phi_ldon_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_ldon_mdz ;
		phi_ldon_mdz:long_name = "phi_ldon_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_ldon_smz ;
		phi_ldon_smz:long_name = "phi_ldon_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_ldon_vir ;
		phi_ldon_vir:long_name = "phi_ldon_vir: Partitioning of viral losses to various dissolved pools" ;
	double phi_ldop_lgz ;
		phi_ldop_lgz:long_name = "phi_ldop_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_ldop_mdz ;
		phi_ldop_mdz:long_name = "phi_ldop_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_ldop_smz ;
		phi_ldop_smz:long_name = "phi_ldop_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_ldop_vir ;
		phi_ldop_vir:long_name = "phi_ldop_vir: Partitioning of viral losses to various dissolved pools" ;
	double phi_lith ;
		phi_lith:long_name = "phi_lith: Remineralization" ;
	double phi_nh4_lgz ;
		phi_nh4_lgz:long_name = "phi_nh4_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_nh4_mdz ;
		phi_nh4_mdz:long_name = "phi_nh4_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_nh4_smz ;
		phi_nh4_smz:long_name = "phi_nh4_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_po4_lgz ;
		phi_po4_lgz:long_name = "phi_po4_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_po4_mdz ;
		phi_po4_mdz:long_name = "phi_po4_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_po4_smz ;
		phi_po4_smz:long_name = "phi_po4_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_sldon_lgz ;
		phi_sldon_lgz:long_name = "phi_sldon_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_sldon_mdz ;
		phi_sldon_mdz:long_name = "phi_sldon_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_sldon_smz ;
		phi_sldon_smz:long_name = "phi_sldon_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_sldon_vir ;
		phi_sldon_vir:long_name = "phi_sldon_vir: Partitioning of viral losses to various dissolved pools" ;
	double phi_sldop_lgz ;
		phi_sldop_lgz:long_name = "phi_sldop_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_sldop_mdz ;
		phi_sldop_mdz:long_name = "phi_sldop_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_sldop_smz ;
		phi_sldop_smz:long_name = "phi_sldop_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_sldop_vir ;
		phi_sldop_vir:long_name = "phi_sldop_vir: Partitioning of viral losses to various dissolved pools" ;
	double phi_srdon_lgz ;
		phi_srdon_lgz:long_name = "phi_srdon_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_srdon_mdz ;
		phi_srdon_mdz:long_name = "phi_srdon_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_srdon_smz ;
		phi_srdon_smz:long_name = "phi_srdon_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_srdon_vir ;
		phi_srdon_vir:long_name = "phi_srdon_vir: Partitioning of viral losses to various dissolved pools" ;
	double phi_srdop_lgz ;
		phi_srdop_lgz:long_name = "phi_srdop_lgz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_srdop_mdz ;
		phi_srdop_mdz:long_name = "phi_srdop_mdz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_srdop_smz ;
		phi_srdop_smz:long_name = "phi_srdop_smz: Partitioning of zooplankton ingestion to other compartments" ;
	double phi_srdop_vir ;
		phi_srdop_vir:long_name = "phi_srdop_vir: Partitioning of viral losses to various dissolved pools" ;
	float po4(ocean_time, s_rho, eta_rho, xi_rho) ;
		po4:long_name = "Phosphate" ;
		po4:units = "mol/kg" ;
		po4:time = "ocean_time" ;
		po4:grid = "grid" ;
		po4:location = "face" ;
		po4:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		po4:field = "po4, scalar, series" ;
		po4:_FillValue = 1.e+37f ;
	double q_p_2_n_bact ;
		q_p_2_n_bact:long_name = "q_p_2_n_bact: Bacteria Stoichiometry - presently static" ;
	double q_p_2_n_lgz ;
		q_p_2_n_lgz:long_name = "q_p_2_n_lgz: Zooplankton Stoichiometry - presently static" ;
	double q_p_2_n_mdz ;
		q_p_2_n_mdz:long_name = "q_p_2_n_mdz: Zooplankton Stoichiometry - presently static" ;
	double q_p_2_n_smz ;
		q_p_2_n_smz:long_name = "q_p_2_n_smz: Zooplankton Stoichiometry - presently static" ;
	double rdrg ;
		rdrg:long_name = "linear drag coefficient" ;
		rdrg:units = "meter second-1" ;
	double rdrg2 ;
		rdrg2:long_name = "quadratic drag coefficient" ;
	double remin_eff_fedet ;
		remin_eff_fedet:long_name = "remin_eff_fedet: Iron chemistry" ;
	float rho(ocean_time, s_rho, eta_rho, xi_rho) ;
		rho:long_name = "density anomaly" ;
		rho:units = "kilogram meter-3" ;
		rho:time = "ocean_time" ;
		rho:grid = "grid" ;
		rho:location = "face" ;
		rho:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		rho:field = "density, scalar, series" ;
		rho:_FillValue = 1.e+37f ;
	double rho0 ;
		rho0:long_name = "mean density used in Boussinesq approximation" ;
		rho0:units = "kilogram meter-3" ;
	double rpcaco3 ;
		rpcaco3:long_name = "rpcaco3: Remineralization" ;
	double rplith ;
		rplith:long_name = "rplith: Remineralization" ;
	double rpsio2 ;
		rpsio2:long_name = "rpsio2: Remineralization" ;
	float s0mk(ocean_time, eta_rho, xi_rho) ;
		s0mk:long_name = "salinity of molecular sub-layer under ice" ;
		s0mk:time = "ocean_time" ;
		s0mk:grid = "grid" ;
		s0mk:location = "face" ;
		s0mk:coordinates = "lon_rho lat_rho ocean_time" ;
		s0mk:field = "salinity, scalar, series" ;
		s0mk:_FillValue = 1.e+37f ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
		s_rho:positive = "up" ;
		s_rho:standard_name = "ocean_s_coordinate_g1" ;
		s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
		s_rho:field = "s_rho, scalar" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
		s_w:positive = "up" ;
		s_w:standard_name = "ocean_s_coordinate_g1" ;
		s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
		s_w:field = "s_w, scalar" ;
	float salt(ocean_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:time = "ocean_time" ;
		salt:grid = "grid" ;
		salt:location = "face" ;
		salt:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		salt:field = "salinity, scalar, series" ;
		salt:_FillValue = 1.e+37f ;
	double si_2_n_max_Lg ;
		si_2_n_max_Lg:long_name = "si_2_n_max_Lg: Other stoichiometry" ;
	double si_2_n_static_Lg ;
		si_2_n_static_Lg:long_name = "si_2_n_static_Lg: Other stoichiometry" ;
	float sidet(ocean_time, s_rho, eta_rho, xi_rho) ;
		sidet:long_name = "Detrital Silicon" ;
		sidet:units = "mol/kg" ;
		sidet:time = "ocean_time" ;
		sidet:grid = "grid" ;
		sidet:location = "face" ;
		sidet:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		sidet:field = "sidet, scalar, series" ;
		sidet:_FillValue = 1.e+37f ;
	float sig11(ocean_time, eta_rho, xi_rho) ;
		sig11:long_name = "internal ice stress 11 component" ;
		sig11:units = "Newton meter-1" ;
		sig11:time = "ocean_time" ;
		sig11:grid = "grid" ;
		sig11:location = "face" ;
		sig11:coordinates = "lon_rho lat_rho ocean_time" ;
		sig11:field = "ice stress 11, scalar, series" ;
		sig11:_FillValue = 1.e+37f ;
	float sig12(ocean_time, eta_rho, xi_rho) ;
		sig12:long_name = "internal ice stress 12 component" ;
		sig12:units = "Newton meter-1" ;
		sig12:time = "ocean_time" ;
		sig12:grid = "grid" ;
		sig12:location = "face" ;
		sig12:coordinates = "lon_rho lat_rho ocean_time" ;
		sig12:field = "ice stress 12, scalar, series" ;
		sig12:_FillValue = 1.e+37f ;
	float sig22(ocean_time, eta_rho, xi_rho) ;
		sig22:long_name = "internal ice stress 22 component" ;
		sig22:units = "Newton meter-1" ;
		sig22:time = "ocean_time" ;
		sig22:grid = "grid" ;
		sig22:location = "face" ;
		sig22:coordinates = "lon_rho lat_rho ocean_time" ;
		sig22:field = "ice stress 22, scalar, series" ;
		sig22:_FillValue = 1.e+37f ;
	float silg(ocean_time, s_rho, eta_rho, xi_rho) ;
		silg:long_name = "Large Phytoplankton Silicon" ;
		silg:units = "mol/kg" ;
		silg:time = "ocean_time" ;
		silg:grid = "grid" ;
		silg:location = "face" ;
		silg:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		silg:field = "silg, scalar, series" ;
		silg:_FillValue = 1.e+37f ;
	float sio4(ocean_time, s_rho, eta_rho, xi_rho) ;
		sio4:long_name = "Silicate" ;
		sio4:units = "mol/kg" ;
		sio4:time = "ocean_time" ;
		sio4:grid = "grid" ;
		sio4:location = "face" ;
		sio4:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		sio4:field = "sio4, scalar, series" ;
		sio4:_FillValue = 1.e+37f ;
	float sldon(ocean_time, s_rho, eta_rho, xi_rho) ;
		sldon:long_name = "Semilabile DON" ;
		sldon:units = "mol/kg" ;
		sldon:time = "ocean_time" ;
		sldon:grid = "grid" ;
		sldon:location = "face" ;
		sldon:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		sldon:field = "sldon, scalar, series" ;
		sldon:_FillValue = 1.e+37f ;
	double smz_ipa_bact ;
		smz_ipa_bact:long_name = "smz_ipa_bact: Zooplankton switching and prey preference parameters" ;
	double smz_ipa_det ;
		smz_ipa_det:long_name = "smz_ipa_det: Zooplankton switching and prey preference parameters" ;
	double smz_ipa_diaz ;
		smz_ipa_diaz:long_name = "smz_ipa_diaz: Zooplankton switching and prey preference parameters" ;
	double smz_ipa_lgp ;
		smz_ipa_lgp:long_name = "smz_ipa_lgp: Zooplankton switching and prey preference parameters" ;
	double smz_ipa_lgz ;
		smz_ipa_lgz:long_name = "smz_ipa_lgz: Zooplankton switching and prey preference parameters" ;
	double smz_ipa_mdz ;
		smz_ipa_mdz:long_name = "smz_ipa_mdz: Zooplankton switching and prey preference parameters" ;
	double smz_ipa_smp ;
		smz_ipa_smp:long_name = "smz_ipa_smp: Zooplankton switching and prey preference parameters" ;
	double smz_ipa_smz ;
		smz_ipa_smz:long_name = "smz_ipa_smz: Zooplankton switching and prey preference parameters" ;
	float snow_thick(ocean_time, eta_rho, xi_rho) ;
		snow_thick:long_name = "thickness of snow cover" ;
		snow_thick:units = "meter" ;
		snow_thick:time = "ocean_time" ;
		snow_thick:grid = "grid" ;
		snow_thick:location = "face" ;
		snow_thick:coordinates = "lon_rho lat_rho ocean_time" ;
		snow_thick:field = "snow thickness, scalar, series" ;
		snow_thick:_FillValue = 1.e+37f ;
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = 0, 1 ;
		spherical:flag_meanings = "Cartesian spherical" ;
	float srdon(ocean_time, s_rho, eta_rho, xi_rho) ;
		srdon:long_name = "Semi-Refractory DON" ;
		srdon:units = "mol/kg" ;
		srdon:time = "ocean_time" ;
		srdon:grid = "grid" ;
		srdon:location = "face" ;
		srdon:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		srdon:field = "srdon, scalar, series" ;
		srdon:_FillValue = 1.e+37f ;
	float t0mk(ocean_time, eta_rho, xi_rho) ;
		t0mk:long_name = "temperature of molecular sub-layer under ice" ;
		t0mk:units = "degrees Celsius" ;
		t0mk:time = "ocean_time" ;
		t0mk:grid = "grid" ;
		t0mk:location = "face" ;
		t0mk:coordinates = "lon_rho lat_rho ocean_time" ;
		t0mk:field = "temperature, scalar, series" ;
		t0mk:_FillValue = 1.e+37f ;
	float tau_iw(ocean_time, eta_rho, xi_rho) ;
		tau_iw:long_name = "ice-water friction velocity" ;
		tau_iw:units = "meter second-1" ;
		tau_iw:time = "ocean_time" ;
		tau_iw:grid = "grid" ;
		tau_iw:location = "face" ;
		tau_iw:coordinates = "lon_rho lat_rho ocean_time" ;
		tau_iw:field = "friction velocity, scalar, series" ;
		tau_iw:_FillValue = 1.e+37f ;
	float temp(ocean_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:time = "ocean_time" ;
		temp:grid = "grid" ;
		temp:location = "face" ;
		temp:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		temp:field = "temperature, scalar, series" ;
		temp:_FillValue = 1.e+37f ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	double thetamax_Di ;
		thetamax_Di:long_name = "thetamax_Di: Phytoplankton light limitation/growth rate" ;
	double thetamax_Lg ;
		thetamax_Lg:long_name = "thetamax_Lg: Phytoplankton light limitation/growth rate" ;
	double thetamax_Sm ;
		thetamax_Sm:long_name = "thetamax_Sm: Phytoplankton light limitation/growth rate" ;
	double thetamin ;
		thetamin:long_name = "thetamin: Phytoplankton light limitation/growth rate" ;
	double thetamin_nolim ;
		thetamin_nolim:long_name = "thetamin_nolim: Phytoplankton light limitation/growth rate" ;
	float ti(ocean_time, eta_rho, xi_rho) ;
		ti:long_name = "interior ice temperature" ;
		ti:units = "degrees Celcius" ;
		ti:time = "ocean_time" ;
		ti:grid = "grid" ;
		ti:location = "face" ;
		ti:coordinates = "lon_rho lat_rho ocean_time" ;
		ti:field = "interior temperature, scalar, series" ;
		ti:_FillValue = 1.e+37f ;
	float tisrf(ocean_time, eta_rho, xi_rho) ;
		tisrf:long_name = "temperature of ice surface" ;
		tisrf:units = "degrees Celcius" ;
		tisrf:time = "ocean_time" ;
		tisrf:grid = "grid" ;
		tisrf:location = "face" ;
		tisrf:coordinates = "lon_rho lat_rho ocean_time" ;
		tisrf:field = "surface temperature, scalar, series" ;
		tisrf:_FillValue = 1.e+37f ;
	float u(ocean_time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:time = "ocean_time" ;
		u:grid = "grid" ;
		u:location = "edge1" ;
		u:coordinates = "lon_u lat_u s_rho ocean_time" ;
		u:field = "u-velocity, scalar, series" ;
		u:_FillValue = 1.e+37f ;
	float ubar(ocean_time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:time = "ocean_time" ;
		ubar:grid = "grid" ;
		ubar:location = "edge1" ;
		ubar:coordinates = "lon_u lat_u ocean_time" ;
		ubar:field = "ubar-velocity, scalar, series" ;
		ubar:_FillValue = 1.e+37f ;
	float uice(ocean_time, eta_u, xi_u) ;
		uice:long_name = "u-component of ice velocity" ;
		uice:units = "meter second-1" ;
		uice:time = "ocean_time" ;
		uice:grid = "grid" ;
		uice:location = "edge1" ;
		uice:coordinates = "lon_u lat_u ocean_time" ;
		uice:field = "u-component of ice velocity, scalar, series" ;
		uice:_FillValue = 1.e+37f ;
	float v(ocean_time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:time = "ocean_time" ;
		v:grid = "grid" ;
		v:location = "edge2" ;
		v:coordinates = "lon_v lat_v s_rho ocean_time" ;
		v:field = "v-velocity, scalar, series" ;
		v:_FillValue = 1.e+37f ;
	float vbar(ocean_time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:time = "ocean_time" ;
		vbar:grid = "grid" ;
		vbar:location = "edge2" ;
		vbar:coordinates = "lon_v lat_v ocean_time" ;
		vbar:field = "vbar-velocity, scalar, series" ;
		vbar:_FillValue = 1.e+37f ;
	float vice(ocean_time, eta_v, xi_v) ;
		vice:long_name = "v-component of ice velocity" ;
		vice:units = "meter second-1" ;
		vice:time = "ocean_time" ;
		vice:grid = "grid" ;
		vice:location = "edge2" ;
		vice:coordinates = "lon_v lat_v ocean_time" ;
		vice:field = "v-component of ice velocity, scalar, series" ;
		vice:_FillValue = 1.e+37f ;
	double vir_Bact ;
		vir_Bact:long_name = "vir_Bact: Phytoplankton and bacterial losses to viruses" ;
	double vir_Di ;
		vir_Di:long_name = "vir_Di: Phytoplankton and bacterial losses to viruses" ;
	double vir_Lg ;
		vir_Lg:long_name = "vir_Lg: Phytoplankton and bacterial losses to viruses" ;
	double vir_Sm ;
		vir_Sm:long_name = "vir_Sm: Phytoplankton and bacterial losses to viruses" ;
	double wsink ;
		wsink:long_name = "wsink: Sinking velocity of detritus" ;
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	double z_sed ;
		z_sed:long_name = "z_sed: Remineralization" ;
	float zeta(ocean_time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:units = "meter" ;
		zeta:time = "ocean_time" ;
		zeta:grid = "grid" ;
		zeta:location = "face" ;
		zeta:coordinates = "lon_rho lat_rho ocean_time" ;
		zeta:field = "free-surface, scalar, series" ;
		zeta:_FillValue = 1.e+37f ;
	double zpllgr ;
		zpllgr:long_name = "zpllgr: Phytoplankton light limitation/growth rate" ;

// global attributes:
		:file = "bgcmip_cobalt/Out/bgcmip_cobalt_03_rst.nc" ;
		:format = "netCDF-3 64bit offset file" ;
		:Conventions = "CF-1.4, SGRID-0.3" ;
		:type = "ROMS/TOMS restart file" ;
		:title = "Bering Sea 10km Grid" ;
		:var_info = "../bering-Apps/Apps/Bering_BGC_variants/varinfo_cobalt_scaledbry.dat" ;
		:rst_file = "bgcmip_cobalt/Out/bgcmip_cobalt_03_rst.nc" ;
		:his_base = "bgcmip_cobalt/Out/bgcmip_cobalt_his" ;
		:avg_base = "bgcmip_cobalt/Out/bgcmip_cobalt_avg" ;
		:dia_base = "bgcmip_cobalt/Out/bgcmip_cobalt_dia" ;
		:sta_file = "bgcmip_cobalt/Out/bgcmip_cobalt_03_sta.nc" ;
		:grd_file = "../../ROMS_Datasets/grids/AlaskaGrids_Bering10K.nc" ;
		:ini_file = "bgcmip_cobalt/Out/bgcmip_cobalt_02_rst.nc" ;
		:tide_file = "../../ROMS_Datasets/OTPS/tides_OTPS_Bering10K.nc" ;
		:frc_file_01 = "../../ROMS_Datasets/BarrowCO2/atmo_co2_barrow_1970_2020.nc" ;
		:frc_file_02 = "../../ROMS_Datasets/Iron/ESM4_Bering10K_iron_dust_clim.nc" ;
		:frc_file_03 = "../../ROMS_Datasets/salinity/sss.clim.nc" ;
		:frc_file_04 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Pair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Pair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Pair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Pair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Pair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Pair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Pair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Pair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Pair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Pair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Pair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Pair-2020.nc" ;
		:frc_file_05 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Qair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Qair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Qair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Qair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Qair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Qair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Qair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Qair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Qair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Qair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Qair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Qair-2020.nc" ;
		:frc_file_06 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Tair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Tair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Tair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Tair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Tair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Tair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Tair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Tair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Tair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Tair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Tair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Tair-2020.nc" ;
		:frc_file_07 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Uwind-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Uwind-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Uwind-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Uwind-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Uwind-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Uwind-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Uwind-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Uwind-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Uwind-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Uwind-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Uwind-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Uwind-2020.nc" ;
		:frc_file_08 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Vwind-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Vwind-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Vwind-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Vwind-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Vwind-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Vwind-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Vwind-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Vwind-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Vwind-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Vwind-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Vwind-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Vwind-2020.nc" ;
		:frc_file_09 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-rain-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-rain-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-rain-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-rain-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-rain-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-rain-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-rain-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-rain-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-rain-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-rain-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-rain-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-rain-2020.nc" ;
		:frc_file_10 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-swrad-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-swrad-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-swrad-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-swrad-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-swrad-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-swrad-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-swrad-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-swrad-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-swrad-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-swrad-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-swrad-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-swrad-2020.nc" ;
		:frc_file_11 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-lwrad-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-lwrad-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-lwrad-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-lwrad-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-lwrad-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-lwrad-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-lwrad-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-lwrad-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-lwrad-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-lwrad-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-lwrad-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-lwrad-2020.nc" ;
		:frc_file_12 = "../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2009.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2010.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2011.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2012.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2013.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2014.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2015.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2016.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2017.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2018.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2019.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2020.nc" ;
		:frc_file_13 = "../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2009.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2010.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2011.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2012.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2013.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2014.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2015.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2016.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2017.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2018.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2019.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2020.nc" ;
		:bry_file_01 = "../../ROMS_Datasets/WOA2018/WOA2018_Bering10K_N30_brybgc.nc" ;
		:bry_file_02 = "../../ROMS_Datasets/CFS/2009/CFS-ocean-Bering10K-N30-bryocn-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-ocean-Bering10K-N30-bryocn-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-ocean-Bering10K-N30-bryocn-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-ocean-Bering10K-N30-bryocn-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-ocean-Bering10K-N30-bryocn-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-ocean-Bering10K-N30-bryocn-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-ocean-Bering10K-N30-bryocn-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-ocean-Bering10K-N30-bryocn-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-ocean-Bering10K-N30-bryocn-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-ocean-Bering10K-N30-bryocn-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-ocean-Bering10K-N30-bryocn-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-ocean-Bering10K-N30-bryocn-2020.nc" ;
		:bry_file_03 = "../../ROMS_Datasets/CFS/2009/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2020.nc" ;
		:clm_file_01 = "../../ROMS_Datasets/initial/ini_hindcast_unnested_Bering10K_BIO_COBALT.nc" ;
		:script_file = "bgcmip_cobalt/In/bgcmip_cobalt_03_ocean.in" ;
		:bpar_file = "bgcmip_cobalt/In/bgcmip_cobalt_bpar.in" ;
		:spos_file = "bgcmip_cobalt/In/bgcmip_cobalt_spos.in" ;
		:NLM_TADV = "\n",
			"ADVECTION:   HORIZONTAL   VERTICAL     \n",
			"temp:        Centered4    Centered4    \n",
			"salt:        Centered4    Centered4    \n",
			"nsm:         HSIMT        HSIMT        \n",
			"nlg:         HSIMT        HSIMT        \n",
			"ndi:         HSIMT        HSIMT        \n",
			"nsmz:        HSIMT        HSIMT        \n",
			"nmdz:        HSIMT        HSIMT        \n",
			"nlgz:        HSIMT        HSIMT        \n",
			"ldon:        HSIMT        HSIMT        \n",
			"sldon:       HSIMT        HSIMT        \n",
			"srdon:       HSIMT        HSIMT        \n",
			"nbact:       HSIMT        HSIMT        \n",
			"nh4:         HSIMT        HSIMT        \n",
			"no3:         HSIMT        HSIMT        \n",
			"ndet:        HSIMT        HSIMT        \n",
			"sio4:        HSIMT        HSIMT        \n",
			"silg:        HSIMT        HSIMT        \n",
			"sidet:       HSIMT        HSIMT        \n",
			"cadet_calc:  HSIMT        HSIMT        \n",
			"cadet_arag:  HSIMT        HSIMT        \n",
			"lith:        HSIMT        HSIMT        \n",
			"lithdet:     HSIMT        HSIMT        \n",
			"po4:         HSIMT        HSIMT        \n",
			"fesm:        HSIMT        HSIMT        \n",
			"fedi:        HSIMT        HSIMT        \n",
			"felg:        HSIMT        HSIMT        \n",
			"fed:         HSIMT        HSIMT        \n",
			"fedet:       HSIMT        HSIMT        \n",
			"o2:          HSIMT        HSIMT        \n",
			"dic:         HSIMT        HSIMT        \n",
			"alk:         HSIMT        HSIMT" ;
		:NLM_LBC = "\n",
			"EDGE:        WEST   SOUTH  EAST   NORTH  \n",
			"zeta:        Che    Che    Clo    Clo    \n",
			"ubar:        Fla    Fla    Clo    Clo    \n",
			"vbar:        Fla    Fla    Clo    Clo    \n",
			"u:           RadNud RadNud Clo    Clo    \n",
			"v:           RadNud RadNud Clo    Clo    \n",
			"temp:        RadNud RadNud Clo    Clo    \n",
			"salt:        RadNud RadNud Clo    Clo    \n",
			"nsm:         RadNud RadNud Clo    Clo    \n",
			"nlg:         RadNud RadNud Clo    Clo    \n",
			"ndi:         RadNud RadNud Clo    Clo    \n",
			"nsmz:        RadNud RadNud Clo    Clo    \n",
			"nmdz:        RadNud RadNud Clo    Clo    \n",
			"nlgz:        RadNud RadNud Clo    Clo    \n",
			"ldon:        RadNud RadNud Clo    Clo    \n",
			"sldon:       RadNud RadNud Clo    Clo    \n",
			"srdon:       RadNud RadNud Clo    Clo    \n",
			"nbact:       RadNud RadNud Clo    Clo    \n",
			"nh4:         RadNud RadNud Clo    Clo    \n",
			"no3:         RadNud RadNud Clo    Clo    \n",
			"ndet:        RadNud RadNud Clo    Clo    \n",
			"sio4:        RadNud RadNud Clo    Clo    \n",
			"silg:        RadNud RadNud Clo    Clo    \n",
			"sidet:       RadNud RadNud Clo    Clo    \n",
			"cadet_calc:  RadNud RadNud Clo    Clo    \n",
			"cadet_arag:  RadNud RadNud Clo    Clo    \n",
			"lith:        RadNud RadNud Clo    Clo    \n",
			"lithdet:     RadNud RadNud Clo    Clo    \n",
			"po4:         RadNud RadNud Clo    Clo    \n",
			"fesm:        RadNud RadNud Clo    Clo    \n",
			"fedi:        RadNud RadNud Clo    Clo    \n",
			"felg:        RadNud RadNud Clo    Clo    \n",
			"fed:         RadNud RadNud Clo    Clo    \n",
			"fedet:       RadNud RadNud Clo    Clo    \n",
			"o2:          RadNud RadNud Clo    Clo    \n",
			"dic:         RadNud RadNud Clo    Clo    \n",
			"alk:         RadNud RadNud Clo    Clo    \n",
			"uice:        Gra    Gra    Clo    Clo    \n",
			"vice:        Gra    Gra    Clo    Clo    \n",
			"aice:        Clo    Clo    Clo    Clo    \n",
			"hice:        Clo    Clo    Clo    Clo    \n",
			"tisrf:       Clo    Clo    Clo    Clo    \n",
			"snow_thick:  Clo    Clo    Clo    Clo    \n",
			"sig11:       Clo    Clo    Clo    Clo    \n",
			"sig12:       Clo    Clo    Clo    Clo    \n",
			"sig22:       Clo    Clo    Clo    Clo" ;
		:git_url = "git@github.com:beringnpz/roms.git" ;
		:git_rev = "cobalttweaks commit c26d625ca5e83a0070032b5ad50faeeec0874813" ;
		:code_dir = "/gscratch/bumblereem/kearney/roms-kate-ice" ;
		:header_dir = "/gscratch/bumblereem/kearney/BGC_hindcasts_workdir" ;
		:header_file = "bering_10k.h" ;
		:os = "Linux" ;
		:cpu = "x86_64" ;
		:compiler_system = "ifort" ;
		:compiler_command = "/gscratch/sw/intel-201703/compilers_and_libraries_2017.2.174/linux/mpi/intel64/b" ;
		:compiler_flags = "-fp-model precise -heap-arrays -ip -O3 -traceback -check uninit -ip -O3" ;
		:tiling = "007x020" ;
		:history = "Fri Sep 22 11:02:56 2023: ncks -F -d ocean_time,1,1 /gscratch/bumblereem/kearney/BGC_hindcasts_workdir/bgcmip_cobalt/Out/bgcmip_cobalt_03_rst.nc ../ini_hindcastloop2_BIO_COBALT.nc\n",
			"ROMS/TOMS, Version 3.9, Tuesday - June 27, 2023 -  2:10:17 AM" ;
		:ana_file = "ROMS/Functionals/ana_btflux.h, /gscratch/bumblereem/kearney/BGC_hindcasts_workdir/ana_psource.h, ROMS/Functionals/ana_srflux.h, ROMS/Functionals/ana_stflux.h, ROMS/Functionals/ana_aiobc.h, ROMS/Functionals/ana_hiobc.h, ROMS/Functionals/ana_hsnobc.h" ;
		:bio_file = "--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------" ;
		:CPP_options = "BERING_10K, ADD_FSOBC, ADD_M2OBC, ALBEDO_CURVE, ANA_BPFLUX, ANA_BSFLUX, ANA_BTFLUX, ANA_PSOURCE, ANA_SPFLUX, ASSUMED_SHAPE, AVERAGES, BIO_COBALT, !BOUNDARY_ALLGATHER, BULK_FLUXES, CCSM_FLUXES, COBALT_CARBON, COBALT_IRON, NO_IRON_COAST, COBALT_MINERALS, COLLECT_ALLGATHER, COASTAL_ATTEN, CORE_FORCING, CURVGRID, DIAGNOSTICS_BIO, DIAGNOSTICS_TS, DIFF_GRID, DIURNAL_SRFLUX, DJ_GRADPS, DOUBLE_PRECISION, EMINUSP, ICE_ADVECT, ICE_BULK_FLUXES, ICE_EVP, ICE_MK, ICE_MODEL, ICE_MOMENTUM, ICE_SMOLAR, ICE_THERMO, LIMIT_BSTRESS, LMD_CONVEC, LMD_MIXING, LMD_NONLOCAL, LMD_RIMIX, LMD_SHAPIRO, LMD_SKPP, LONGWAVE_OUT, MASKING, MIX_GEO_TS, MIX_S_UV, MPI, NONLINEAR, NONLIN_EOS, NO_WRITE_GRID, OPTIC_MANIZZA, POT_TIDES, POWER_LAW, PROFILE, RADIATION_2D, REDUCE_ALLGATHER, RUNOFF, RST_SINGLE, SALINITY, SCORRECTION, SOLAR_SOURCE, SOLVE3D, SSH_TIDES, STATIONS, TIDES_ASTRO, TS_DIF2, UV_ADV, UV_COR, UV_U3HADVECTION, UV_SADVECTION, UV_DRAG_GRID, UV_LDRAG, UV_TIDES, UV_VIS2, UV_SMAGORINSKY, VAR_RHO_2D, VISC_GRID, VISC_3DCOEF" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
