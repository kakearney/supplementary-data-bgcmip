netcdf CFS-atmos-northPacific-Uwind-2017 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:missing_value = -1.e+34 ;
		Uwind:_FillValue = -1.e+34 ;
		Uwind:time = "wind_time" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:height_above_ground1 = 10.f ;
		Uwind:long_name = "U wind" ;
		Uwind:history = "From roms-cfs-atmos-Uwind-2017" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:10:08 2022: ncks -F -O -d wind_time,3,1462 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2017/roms-cfs-atmos-Uwind-2017.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Uwind-2017.nc\n",
			"Mon Sep 17 12:09:49 2018: Time overhang added\n",
			"Mon Sep 17 12:09:42 2018: ncrcat /tmp/tp80e4ff69_3c78_4d3e_8385_b39e2ec684bd.nc frc/roms-cfs-atmos-Uwind-2017.nc /tmp/tp70435bab_9568_48b6_bc64_efc0c77688f4.nc /tmp/tp42b55a5d_c2c9_4940_820d_b4b4be35beaf.nc\n",
			"Mon Sep 17 12:09:41 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2017.nc /tmp/tp80e4ff69_3c78_4d3e_8385_b39e2ec684bd.nc\n",
			"FERRET V7.4  10-Aug-18" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
