netcdf CFS-atmos-northPacific-lwrad-1995 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:38:10 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1995/roms-cfs-atmos-lwrad-1995.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1995/CFS-atmos-northPacific-lwrad-1995.nc\n",
			"Mon Sep 10 13:46:31 2018: Time overhang added\n",
			"Mon Sep 10 13:46:27 2018: ncrcat /tmp/tp073a9574_37e6_4eae_bc3a_b2f2704bd8d1.nc frc/roms-cfs-atmos-lwrad-1995.nc /tmp/tp00c137c7_70ab_4192_9419_92d9dec0b2b4.nc /tmp/tp8d5a0cb3_c3fc_4b65_80b7_e1a301297c3e.nc\n",
			"Mon Sep 10 13:46:27 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-1995.nc /tmp/tp073a9574_37e6_4eae_bc3a_b2f2704bd8d1.nc\n",
			"Thu Sep  6 09:52:39 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1995_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-1995.nc\n",
			"04-Oct-2017 17:37:48: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
