netcdf CFS-atmos-northPacific-lwrad-1997 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:34 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1997/roms-cfs-atmos-lwrad-1997.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1997/CFS-atmos-northPacific-lwrad-1997.nc\n",
			"Mon Sep 10 13:46:43 2018: Time overhang added\n",
			"Mon Sep 10 13:46:39 2018: ncrcat /tmp/tpcd576839_a1f0_4557_ad1a_f622d635b1bd.nc frc/roms-cfs-atmos-lwrad-1997.nc /tmp/tp9ced36ae_385f_4aad_b31d_883d25e0942a.nc /tmp/tp835e46c8_1ba6_40a7_b0ac_9dc3264d1205.nc\n",
			"Mon Sep 10 13:46:39 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-1997.nc /tmp/tpcd576839_a1f0_4557_ad1a_f622d635b1bd.nc\n",
			"Thu Sep  6 10:09:42 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1997_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-1997.nc\n",
			"04-Oct-2017 17:42:40: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
