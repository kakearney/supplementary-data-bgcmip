netcdf CFS-ocean-ESPER-NEP-N30-brycarbon-2014 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 642 ;
	xi_rho = 226 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 16:28:22 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 16:25:26 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2014/CFS-ocean-NEP-N30-bryocn-2014.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2014/CFS-ocean-ESPER-NEP-N30-brycarbon-2014.nc\n",
			"Mon Jan  9 10:12:24 2023: ncrcat -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad02.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad03.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad04.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad05.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad06.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad07.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad08.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad09.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad10.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad11.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad12.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad13.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad14.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad15.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad16.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad17.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad18.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad19.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad20.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad21.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad22.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad23.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad24.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad25.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad26.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad27.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad28.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad29.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad30.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad31.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad32.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad33.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad34.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad35.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad36.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad37.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad38.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad39.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad40.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad41.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad42.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad43.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad44.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad45.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad46.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad47.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad48.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad49.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad50.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad51.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad52.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad53.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad54.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad55.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad56.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad57.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad58.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad59.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad60.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad61.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad62.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad63.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad64.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad65.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad66.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad67.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad68.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad69.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad70.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad71.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad72.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad73.nc <>/final/2014/CFS-ocean-NEP-N30-bryocn-2014.nc\n",
			"Mon Jan  9 10:09:48 2023: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad01.nc\n",
			"Mon Jan  9 10:09:46 2023: ncra -O <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad01.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad01.nc\n",
			"Mon Jan  9 10:09:45 2023: ncrcat -O <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010100.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010106.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010112.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010118.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010200.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010206.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010212.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010218.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010300.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010306.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010312.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010318.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010400.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010406.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010412.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010418.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010500.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010506.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010512.nc <>/prep/singletime/CFS-ocean-NEP-N30-bryocn-2014010518.nc <>/prep/pentads/CFS-ocean-NEP-N30-bryocn-2014pentad01.nc\n",
			"Sun Jan 08 19:52:54 2023: CFS data added\n",
			"Tue Dec 20 15:09:10 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
