netcdf CFS-atmos-northPacific-Qair-1994 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:missing_value = -1.e+34 ;
		Qair:_FillValue = -1.e+34 ;
		Qair:time = "qair_time" ;
		Qair:coordinates = "lon lat" ;
		Qair:height_above_ground = 2.f ;
		Qair:long_name = "specific humidity" ;
		Qair:history = "From roms-cfs-atmos-Qair-1994" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double qair_time(qair_time) ;
		qair_time:units = "day since 1900-01-01 00:00:00" ;
		qair_time:time_origin = "01-JAN-1900 00:00:00" ;
		qair_time:axis = "T" ;
		qair_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:34:44 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1994/roms-cfs-atmos-Qair-1994.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1994/CFS-atmos-northPacific-Qair-1994.nc\n",
			"Wed Nov 20 14:04:52 2019: Time overhang added to both ends\n",
			"Wed Nov 20 14:04:47 2019: ncrcat /tmp/tpc74673a6_0d81_476d_9351_694d077c9430.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1994/roms-cfs-atmos-Qair-1994.nc /tmp/tp9ccdac28_dbdb_447e_8deb_61cede0c14c0.nc /tmp/tp1b03f26a_a617_4725_9658_cbb4d33b5514.nc\n",
			"Wed Nov 20 14:04:45 2019: ncks -F -d qair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1994/roms-cfs-atmos-Qair-1994.nc /tmp/tpc74673a6_0d81_476d_9351_694d077c9430.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
