netcdf CFS-atmos-northPacific-Tair-2004 {
dimensions:
	tair_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:50:47 2022: ncks -F -O -d tair_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2004/roms-cfs-atmos-Tair-2004.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2004/CFS-atmos-northPacific-Tair-2004.nc\n",
			"Mon Sep 10 13:38:17 2018: Time overhang added\n",
			"Mon Sep 10 13:38:14 2018: ncrcat /tmp/tpb0f1a7b5_ed35_4319_8ba1_bcc288a86761.nc frc/roms-cfs-atmos-Tair-2004.nc /tmp/tp9f697700_d169_4296_a37a_57e85cc7d7f6.nc /tmp/tpb386dde5_adc9_467f_90de_332d866a1af8.nc\n",
			"Mon Sep 10 13:38:13 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2004.nc /tmp/tpb0f1a7b5_ed35_4319_8ba1_bcc288a86761.nc\n",
			"Thu Sep  6 11:10:14 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2004.nc\n",
			"Thu Sep  6 11:09:20 2018: ncks -O -F -d air_time,2,1465 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2004_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2004.nc\n",
			"04-Oct-2017 17:59:35: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
