netcdf CFS-atmos-northPacific-Pair-1997 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:00 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1997/roms-cfs-atmos-Pair-1997.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1997/CFS-atmos-northPacific-Pair-1997.nc\n",
			"Mon Sep 10 13:31:43 2018: Time overhang added\n",
			"Mon Sep 10 13:31:38 2018: ncrcat /tmp/tp74b30236_a479_4112_b269_d1f09cedec8b.nc frc/roms-cfs-atmos-Pair-1997.nc /tmp/tp96c2fbea_f6eb_4175_a289_6aa8f072bb47.nc /tmp/tp6ae71bd3_2e11_4184_8e48_a8e345d281e7.nc\n",
			"Mon Sep 10 13:31:38 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-1997.nc /tmp/tp74b30236_a479_4112_b269_d1f09cedec8b.nc\n",
			"Thu Sep  6 10:06:34 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1997.nc\n",
			"Thu Sep  6 10:05:30 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1997_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1997.nc\n",
			"04-Oct-2017 17:41:45: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
