netcdf CFS-atmos-northPacific-Pair-2009 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:58:00 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2009/roms-cfs-atmos-Pair-2009.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Pair-2009.nc\n",
			"Mon Sep 10 13:32:54 2018: Time overhang added\n",
			"Mon Sep 10 13:32:51 2018: ncrcat /tmp/tpe505c5ae_946d_492e_b680_ba82dac3ea8f.nc frc/roms-cfs-atmos-Pair-2009.nc /tmp/tpd357b1f2_b06a_49f9_a725_064481332c68.nc /tmp/tpad0ee0ac_23a3_4f1e_9f46_741e855752ea.nc\n",
			"Mon Sep 10 13:32:50 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2009.nc /tmp/tpe505c5ae_946d_492e_b680_ba82dac3ea8f.nc\n",
			"Thu Sep  6 11:58:31 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2009.nc\n",
			"Thu Sep  6 11:57:32 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2009_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2009.nc\n",
			"04-Oct-2017 18:09:27: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
