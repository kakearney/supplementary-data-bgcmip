netcdf CFS-atmos-northPacific-Vwind-1995 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:37:23 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1995/roms-cfs-atmos-Vwind-1995.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1995/CFS-atmos-northPacific-Vwind-1995.nc\n",
			"Mon Sep 10 13:43:27 2018: Time overhang added\n",
			"Mon Sep 10 13:43:23 2018: ncrcat /tmp/tpae931693_94cc_4ec4_af87_db5c84cf924e.nc frc/roms-cfs-atmos-Vwind-1995.nc /tmp/tpa226b156_4045_41ad_818c_7024bdf143f1.nc /tmp/tpcc1f9cdd_8382_4a69_89dc_a30d23bf22cd.nc\n",
			"Mon Sep 10 13:43:23 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-1995.nc /tmp/tpae931693_94cc_4ec4_af87_db5c84cf924e.nc\n",
			"Thu Sep  6 09:54:56 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1995_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-1995.nc\n",
			"04-Oct-2017 17:38:16: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
