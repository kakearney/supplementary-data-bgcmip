netcdf CFS-atmos-northPacific-Vwind-2008 {
dimensions:
	wind_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:57:07 2022: ncks -F -O -d wind_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2008/roms-cfs-atmos-Vwind-2008.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2008/CFS-atmos-northPacific-Vwind-2008.nc\n",
			"Mon Sep 10 13:44:41 2018: Time overhang added\n",
			"Mon Sep 10 13:44:38 2018: ncrcat /tmp/tp6b0e68a7_1a86_48d7_bc35_432d84df688c.nc frc/roms-cfs-atmos-Vwind-2008.nc /tmp/tp4bce1d4b_2a17_4f9f_a812_1b7823f1fbd9.nc /tmp/tp800f07dc_55d4_4bbb_b116_8441b75c774f.nc\n",
			"Mon Sep 10 13:44:37 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2008.nc /tmp/tp6b0e68a7_1a86_48d7_bc35_432d84df688c.nc\n",
			"Thu Sep  6 11:56:39 2018: ncks -O -F -d wind_time,2,1465 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2008_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2008.nc\n",
			"04-Oct-2017 18:08:30: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
