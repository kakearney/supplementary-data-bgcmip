netcdf CFS-atmos-northPacific-Uwind-2020 {
dimensions:
	wind_time = UNLIMITED ; // (1448 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:missing_value = -1.e+34 ;
		Uwind:_FillValue = -1.e+34 ;
		Uwind:time = "wind_time" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:height_above_ground1 = 10.f ;
		Uwind:long_name = "U wind" ;
		Uwind:history = "From roms-cfs-atmos-Uwind-2020" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:54:37 2022: ncks -F -O -d wind_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Uwind-2020.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Uwind-2020.nc\n",
			"Wed Jan 27 10:11:34 2021: Time overhang added to both ends\n",
			"Wed Jan 27 10:11:25 2021: ncrcat /tmp/tp4ecda692_4b24_4080_ae4f_24e5a253c1c0.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Uwind-2020.nc /tmp/tpe70de67c_c014_4f23_8fa9_088d7a40e196.nc /tmp/tp42724d90_13f8_42c3_9cd6_107e8d6cb187.nc\n",
			"Wed Jan 27 10:11:24 2021: ncks -F -d wind_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Uwind-2020.nc /tmp/tp4ecda692_4b24_4080_ae4f_24e5a253c1c0.nc\n",
			"FERRET V7.6  26-Jan-21" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
