netcdf CFS-atmos-northPacific-Qair-2016 {
dimensions:
	qair_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Mon Oct 31 11:54:09 2022: ncks -F -O -d qair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2016/roms-cfs-atmos-Qair-2016.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Qair-2016.nc\n",
			"Mon Sep 10 13:37:01 2018: Time overhang added\n",
			"Mon Sep 10 13:36:53 2018: ncrcat /tmp/tp6bd6ab6d_1667_4ce1_afc2_20543df0cba9.nc frc/roms-cfs-atmos-Qair-2016.nc /tmp/tp60e51f9b_e13d_4bc8_a880_cef689faa4f5.nc /tmp/tp9c01323f_ca20_4f6f_b485_3011ef06ab26.nc\n",
			"Mon Sep 10 13:36:53 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2016.nc /tmp/tp6bd6ab6d_1667_4ce1_afc2_20543df0cba9.nc\n",
			"Thu Sep  6 14:11:27 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2016.nc\n",
			"Thu Sep  6 14:09:32 2018: ncks -O -F -d air_time,2,1449 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2016_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2016.nc\n",
			"04-Oct-2017 18:32:42: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
