netcdf ini_hindcastloop2_BIO_BANAS {
dimensions:
	ocean_time = UNLIMITED ; // (1 currently)
	s_w = 31 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
	tracer = 8 ;
	s_rho = 30 ;
	boundary = 4 ;
	eta_u = 258 ;
	xi_u = 181 ;
	eta_v = 257 ;
	xi_v = 182 ;
variables:
	float AKs(ocean_time, s_w, eta_rho, xi_rho) ;
		AKs:long_name = "salinity vertical diffusion coefficient" ;
		AKs:units = "meter2 second-1" ;
		AKs:time = "ocean_time" ;
		AKs:grid = "grid" ;
		AKs:location = "face" ;
		AKs:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKs:field = "AKs, scalar, series" ;
	float AKt(ocean_time, s_w, eta_rho, xi_rho) ;
		AKt:long_name = "temperature vertical diffusion coefficient" ;
		AKt:units = "meter2 second-1" ;
		AKt:time = "ocean_time" ;
		AKt:grid = "grid" ;
		AKt:location = "face" ;
		AKt:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKt:field = "AKt, scalar, series" ;
	float AKv(ocean_time, s_w, eta_rho, xi_rho) ;
		AKv:long_name = "vertical viscosity coefficient" ;
		AKv:units = "meter2 second-1" ;
		AKv:time = "ocean_time" ;
		AKv:grid = "grid" ;
		AKv:location = "face" ;
		AKv:coordinates = "lon_rho lat_rho s_w ocean_time" ;
		AKv:field = "AKv, scalar, series" ;
	double Akt_bak(tracer) ;
		Akt_bak:long_name = "background vertical mixing coefficient for tracers" ;
		Akt_bak:units = "meter2 second-1" ;
	double Akv_bak ;
		Akv_bak:long_name = "background vertical mixing coefficient for momentum" ;
		Akv_bak:units = "meter2 second-1" ;
	int BioIter ;
		BioIter:long_name = "number of iterations to achieve convergence" ;
	int CNratio ;
		CNratio:long_name = "phytoplankton C:N ratio" ;
		CNratio:units = "molC/molN" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
		Cs_r:field = "Cs_r, scalar" ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
		Cs_w:field = "Cs_w, scalar" ;
	int Ecrit ;
		Ecrit:long_name = "light level of alpha_win/alpha_sum transition" ;
		Ecrit:units = "W m^-2" ;
	double FSobc_in(boundary) ;
		FSobc_in:long_name = "free-surface inflow, nudging inverse time scale" ;
		FSobc_in:units = "second-1" ;
	double FSobc_out(boundary) ;
		FSobc_out:long_name = "free-surface outflow, nudging inverse time scale" ;
		FSobc_out:units = "second-1" ;
	double Falpha ;
		Falpha:long_name = "Power-law shape barotropic filter parameter" ;
	double Fbeta ;
		Fbeta:long_name = "Power-law shape barotropic filter parameter" ;
	double Fgamma ;
		Fgamma:long_name = "Power-law shape barotropic filter parameter" ;
	float Hsbl(ocean_time, eta_rho, xi_rho) ;
		Hsbl:long_name = "depth of oceanic surface boundary layer" ;
		Hsbl:units = "meter" ;
		Hsbl:time = "ocean_time" ;
		Hsbl:grid = "grid" ;
		Hsbl:location = "face" ;
		Hsbl:coordinates = "lon_rho lat_rho ocean_time" ;
		Hsbl:field = "Hsbl, scalar, series" ;
		Hsbl:_FillValue = 1.e+37f ;
	int I0 ;
		I0:long_name = "max microzooplankton ingestion rate" ;
		I0:units = "d^-1" ;
	int Kgraz ;
		Kgraz:long_name = "grazing half-saturation" ;
		Kgraz:units = "uM N" ;
	int Lm2CLM ;
		Lm2CLM:long_name = "2D momentum climatology processing switch" ;
		Lm2CLM:flag_values = 0, 1 ;
		Lm2CLM:flag_meanings = ".FALSE. .TRUE." ;
	int Lm3CLM ;
		Lm3CLM:long_name = "3D momentum climatology processing switch" ;
		Lm3CLM:flag_values = 0, 1 ;
		Lm3CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeM2CLM ;
		LnudgeM2CLM:long_name = "2D momentum climatology nudging activation switch" ;
		LnudgeM2CLM:flag_values = 0, 1 ;
		LnudgeM2CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeM3CLM ;
		LnudgeM3CLM:long_name = "3D momentum climatology nudging activation switch" ;
		LnudgeM3CLM:flag_values = 0, 1 ;
		LnudgeM3CLM:flag_meanings = ".FALSE. .TRUE." ;
	int LnudgeTCLM(tracer) ;
		LnudgeTCLM:long_name = "tracer climatology nudging activation switch" ;
		LnudgeTCLM:flag_values = 0, 1 ;
		LnudgeTCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LsshCLM ;
		LsshCLM:long_name = "sea surface height climatology processing switch" ;
		LsshCLM:flag_values = 0, 1 ;
		LsshCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerCLM(tracer) ;
		LtracerCLM:long_name = "tracer climatology processing switch" ;
		LtracerCLM:flag_values = 0, 1 ;
		LtracerCLM:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerSponge(tracer) ;
		LtracerSponge:long_name = "horizontal diffusivity sponge activation switch" ;
		LtracerSponge:flag_values = 0, 1 ;
		LtracerSponge:flag_meanings = ".FALSE. .TRUE." ;
	int LtracerSrc(tracer) ;
		LtracerSrc:long_name = "tracer point sources and sink activation switch" ;
		LtracerSrc:flag_values = 0, 1 ;
		LtracerSrc:flag_meanings = ".FALSE. .TRUE." ;
	int LuvSponge ;
		LuvSponge:long_name = "horizontal viscosity sponge activation switch" ;
		LuvSponge:flag_values = 0, 1 ;
		LuvSponge:flag_meanings = ".FALSE. .TRUE." ;
	int LuvSrc ;
		LuvSrc:long_name = "momentum point sources and sink activation switch" ;
		LuvSrc:flag_values = 0, 1 ;
		LuvSrc:flag_meanings = ".FALSE. .TRUE." ;
	int LwSrc ;
		LwSrc:long_name = "mass point sources and sink activation switch" ;
		LwSrc:flag_values = 0, 1 ;
		LwSrc:flag_meanings = ".FALSE. .TRUE." ;
	double M2nudg ;
		M2nudg:long_name = "2D momentum nudging/relaxation inverse time scale" ;
		M2nudg:units = "day-1" ;
	double M2obc_in(boundary) ;
		M2obc_in:long_name = "2D momentum inflow, nudging inverse time scale" ;
		M2obc_in:units = "second-1" ;
	double M2obc_out(boundary) ;
		M2obc_out:long_name = "2D momentum outflow, nudging inverse time scale" ;
		M2obc_out:units = "second-1" ;
	double M3nudg ;
		M3nudg:long_name = "3D momentum nudging/relaxation inverse time scale" ;
		M3nudg:units = "day-1" ;
	double M3obc_in(boundary) ;
		M3obc_in:long_name = "3D momentum inflow, nudging inverse time scale" ;
		M3obc_in:units = "second-1" ;
	double M3obc_out(boundary) ;
		M3obc_out:long_name = "3D momentum outflow, nudging inverse time scale" ;
		M3obc_out:units = "second-1" ;
	float NH4(ocean_time, s_rho, eta_rho, xi_rho) ;
		NH4:long_name = "ammonium" ;
		NH4:units = "mmol N m^-3" ;
		NH4:time = "ocean_time" ;
		NH4:grid = "grid" ;
		NH4:location = "face" ;
		NH4:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		NH4:field = "ammonium" ;
		NH4:_FillValue = 1.e+37f ;
	float NO3(ocean_time, s_rho, eta_rho, xi_rho) ;
		NO3:long_name = "nitrate" ;
		NO3:units = "mmol N m^-3" ;
		NO3:time = "ocean_time" ;
		NO3:grid = "grid" ;
		NO3:location = "face" ;
		NO3:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		NO3:field = "nitrate" ;
		NO3:_FillValue = 1.e+37f ;
	int Q_P ;
		Q_P:long_name = "Q10 for phytoplankton" ;
		Q_P:units = "unitless" ;
	int Q_R ;
		Q_R:long_name = "Q10 for bacterial respiration" ;
		Q_R:units = "unitless" ;
	int Q_Z ;
		Q_Z:long_name = "Q10 for zooplankton" ;
		Q_Z:units = "unitless" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double Tnudg(tracer) ;
		Tnudg:long_name = "Tracers nudging/relaxation inverse time scale" ;
		Tnudg:units = "day-1" ;
	double Tnudg_SSS ;
		Tnudg_SSS:long_name = "SSS nudging/relaxation inverse time scale" ;
		Tnudg_SSS:units = "day-1" ;
	double Tobc_in(boundary, tracer) ;
		Tobc_in:long_name = "tracers inflow, nudging inverse time scale" ;
		Tobc_in:units = "second-1" ;
	double Tobc_out(boundary, tracer) ;
		Tobc_out:long_name = "tracers outflow, nudging inverse time scale" ;
		Tobc_out:units = "second-1" ;
	int Vstretching ;
		Vstretching:long_name = "vertical terrain-following stretching function" ;
	int Vtransform ;
		Vtransform:long_name = "vertical terrain-following transformation equation" ;
	double Znudg ;
		Znudg:long_name = "free-surface nudging/relaxation inverse time scale" ;
		Znudg:units = "day-1" ;
	double Zob ;
		Zob:long_name = "bottom roughness" ;
		Zob:units = "meter" ;
	double Zos ;
		Zos:long_name = "surface roughness" ;
		Zos:units = "meter" ;
	float ageice(ocean_time, eta_rho, xi_rho) ;
		ageice:long_name = "age of the ice" ;
		ageice:units = "sec" ;
		ageice:time = "ocean_time" ;
		ageice:grid = "grid" ;
		ageice:location = "face" ;
		ageice:coordinates = "lon_rho lat_rho ocean_time" ;
		ageice:field = "ice age, scalar, series" ;
		ageice:_FillValue = 1.e+37f ;
	float aice(ocean_time, eta_rho, xi_rho) ;
		aice:long_name = "fraction of cell covered by ice" ;
		aice:time = "ocean_time" ;
		aice:grid = "grid" ;
		aice:location = "face" ;
		aice:coordinates = "lon_rho lat_rho ocean_time" ;
		aice:field = "ice concentration, scalar, series" ;
		aice:_FillValue = 1.e+37f ;
	int alpha_sum ;
		alpha_sum:long_name = "initial growth-light slope, summer" ;
		alpha_sum:units = "(W M^-2)^-1 d^-1" ;
	int alpha_win ;
		alpha_win:long_name = "initial growth-light slope, winter" ;
		alpha_win:units = "(W M^-2)^-1 d^-1" ;
	int att_p ;
		att_p:long_name = "light attneuation by phytoplankton" ;
		att_p:units = "m^-1 uM N^-1" ;
	int att_sw ;
		att_sw:long_name = "light attenuation by seawater" ;
		att_sw:units = "m^-1" ;
	int chlNratio ;
		chlNratio:long_name = "chlorohpyll:N ratio" ;
		chlNratio:units = "mg chl/uM N" ;
	float chu_iw(ocean_time, eta_rho, xi_rho) ;
		chu_iw:long_name = "ice-water momentum transfer coefficient" ;
		chu_iw:units = "meter second-1" ;
		chu_iw:time = "ocean_time" ;
		chu_iw:grid = "grid" ;
		chu_iw:location = "face" ;
		chu_iw:coordinates = "lon_rho lat_rho ocean_time" ;
		chu_iw:field = "transfer coefficient, scalar, series" ;
		chu_iw:_FillValue = 1.e+37f ;
	int deltaE ;
		deltaE:long_name = "width of alpha_win/alpha_sum transition" ;
		deltaE:units = "W m^-2" ;
	float det_large(ocean_time, s_rho, eta_rho, xi_rho) ;
		det_large:long_name = "large detritus (aggregates)" ;
		det_large:units = "mmol N m^-3" ;
		det_large:time = "ocean_time" ;
		det_large:grid = "grid" ;
		det_large:location = "face" ;
		det_large:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		det_large:field = "large detritus" ;
		det_large:_FillValue = 1.e+37f ;
	float det_small(ocean_time, s_rho, eta_rho, xi_rho) ;
		det_small:long_name = "small detritus" ;
		det_small:units = "mmol N m^-3" ;
		det_small:time = "ocean_time" ;
		det_small:grid = "grid" ;
		det_small:location = "face" ;
		det_small:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		det_small:field = "small detritus" ;
		det_small:_FillValue = 1.e+37f ;
	double dstart ;
		dstart:long_name = "time stamp assigned to model initilization" ;
		dstart:units = "days since 1900-01-01 00:00:00" ;
		dstart:calendar = "proleptic_gregorian" ;
	double dt ;
		dt:long_name = "size of long time-steps" ;
		dt:units = "second" ;
	double dtfast ;
		dtfast:long_name = "size of short time-steps" ;
		dtfast:units = "second" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	int epsil ;
		epsil:long_name = "microzooplankton growth efficiency" ;
		epsil:units = "unitless" ;
	int fex ;
		fex:long_name = "fraction of grazing excreted to NH4" ;
		fex:units = "unitless" ;
	double gamma2 ;
		gamma2:long_name = "slipperiness parameter" ;
	int grid ;
		grid:cf_role = "grid_topology" ;
		grid:topology_dimension = 2 ;
		grid:node_dimensions = "xi_psi eta_psi" ;
		grid:face_dimensions = "xi_rho: xi_psi (padding: both) eta_rho: eta_psi (padding: both)" ;
		grid:edge1_dimensions = "xi_u: xi_psi eta_u: eta_psi (padding: both)" ;
		grid:edge2_dimensions = "xi_v: xi_psi (padding: both) eta_v: eta_psi" ;
		grid:node_coordinates = "lon_psi lat_psi" ;
		grid:face_coordinates = "lon_rho lat_rho" ;
		grid:edge1_coordinates = "lon_u lat_u" ;
		grid:edge2_coordinates = "lon_v lat_v" ;
		grid:vertical_dimensions = "s_rho: s_w (padding: none)" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	float hice(ocean_time, eta_rho, xi_rho) ;
		hice:long_name = "average ice thickness in cell" ;
		hice:units = "meter" ;
		hice:time = "ocean_time" ;
		hice:grid = "grid" ;
		hice:location = "face" ;
		hice:coordinates = "lon_rho lat_rho ocean_time" ;
		hice:field = "ice thickness, scalar, series" ;
		hice:_FillValue = 1.e+37f ;
	double k_sed1 ;
		k_sed1:long_name = "Depth-based attenuation coefficient, factor" ;
		k_sed1:units = "m^-1" ;
	double k_sed2 ;
		k_sed2:long_name = "Depth-based attenuation coefficient, exponent" ;
		k_sed2:units = "unitless" ;
	int kmin ;
		kmin:long_name = "minmimum half-saturation for NO3" ;
		kmin:units = "uM N" ;
	int m_P ;
		m_P:long_name = "phytoplankton mortality" ;
		m_P:units = "d^-1" ;
	int m_Z ;
		m_Z:long_name = "microzooplankton mortality" ;
		m_Z:units = "d^-1" ;
	int m_agg ;
		m_agg:long_name = "phytoplankton loss via aggregation" ;
		m_agg:units = "(uM N)^-1 d^-1" ;
	float microzoo(ocean_time, s_rho, eta_rho, xi_rho) ;
		microzoo:long_name = "microzooplankton" ;
		microzoo:units = "mmol N m^-3" ;
		microzoo:time = "ocean_time" ;
		microzoo:grid = "grid" ;
		microzoo:location = "face" ;
		microzoo:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		microzoo:field = "microzooplankton" ;
		microzoo:_FillValue = 1.e+37f ;
	int mu0 ;
		mu0:long_name = "maximum phytoplankton growth rate" ;
		mu0:units = "d^-1" ;
	int nAVG ;
		nAVG:long_name = "number of time-steps between time-averaged records" ;
	int nDIA ;
		nDIA:long_name = "number of time-steps between diagnostic records" ;
	int nHIS ;
		nHIS:long_name = "number of time-steps between history records" ;
	int nRST ;
		nRST:long_name = "number of time-steps between restart records" ;
		nRST:cycle = "only latest two records are maintained" ;
	int nSTA ;
		nSTA:long_name = "number of time-steps between stations records" ;
	int ndefAVG ;
		ndefAVG:long_name = "number of time-steps between the creation of average files" ;
	int ndefDIA ;
		ndefDIA:long_name = "number of time-steps between the creation of diagnostic files" ;
	int ndefHIS ;
		ndefHIS:long_name = "number of time-steps between the creation of history files" ;
	int ndtfast ;
		ndtfast:long_name = "number of short time-steps" ;
	double nl_tnu2(tracer) ;
		nl_tnu2:long_name = "nonlinear model Laplacian mixing coefficient for tracers" ;
		nl_tnu2:units = "meter2 second-1" ;
	double nl_visc2 ;
		nl_visc2:long_name = "nonlinear model Laplacian mixing coefficient for momentum" ;
		nl_visc2:units = "meter2 second-1" ;
	int ntimes ;
		ntimes:long_name = "number of long time-steps" ;
	int ntsAVG ;
		ntsAVG:long_name = "starting time-step for accumulation of time-averaged fields" ;
	int ntsDIA ;
		ntsDIA:long_name = "starting time-step for accumulation of diagnostic fields" ;
	double ocean_time(ocean_time) ;
		ocean_time:long_name = "time since initialization" ;
		ocean_time:units = "seconds since 1900-01-01 00:00:00" ;
		ocean_time:calendar = "proleptic_gregorian" ;
		ocean_time:field = "time, scalar, series" ;
	int phi_NH4 ;
		phi_NH4:long_name = "preference for NH4" ;
		phi_NH4:units = "unitless" ;
	float phyto(ocean_time, s_rho, eta_rho, xi_rho) ;
		phyto:long_name = "phytoplankton" ;
		phyto:units = "mmol N m^-3" ;
		phyto:time = "ocean_time" ;
		phyto:grid = "grid" ;
		phyto:location = "face" ;
		phyto:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		phyto:field = "phytoplankton" ;
		phyto:_FillValue = 1.e+37f ;
	int r_nitr ;
		r_nitr:long_name = "nitrification rate" ;
		r_nitr:units = "d^-1" ;
	int r_remin ;
		r_remin:long_name = "detrital remineralization rate" ;
		r_remin:units = "d^-1" ;
	double rdrg ;
		rdrg:long_name = "linear drag coefficient" ;
		rdrg:units = "meter second-1" ;
	double rdrg2 ;
		rdrg2:long_name = "quadratic drag coefficient" ;
	float rho(ocean_time, s_rho, eta_rho, xi_rho) ;
		rho:long_name = "density anomaly" ;
		rho:units = "kilogram meter-3" ;
		rho:time = "ocean_time" ;
		rho:grid = "grid" ;
		rho:location = "face" ;
		rho:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		rho:field = "density, scalar, series" ;
		rho:_FillValue = 1.e+37f ;
	double rho0 ;
		rho0:long_name = "mean density used in Boussinesq approximation" ;
		rho0:units = "kilogram meter-3" ;
	float s0mk(ocean_time, eta_rho, xi_rho) ;
		s0mk:long_name = "salinity of molecular sub-layer under ice" ;
		s0mk:time = "ocean_time" ;
		s0mk:grid = "grid" ;
		s0mk:location = "face" ;
		s0mk:coordinates = "lon_rho lat_rho ocean_time" ;
		s0mk:field = "salinity, scalar, series" ;
		s0mk:_FillValue = 1.e+37f ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
		s_rho:positive = "up" ;
		s_rho:standard_name = "ocean_s_coordinate_g1" ;
		s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
		s_rho:field = "s_rho, scalar" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
		s_w:positive = "up" ;
		s_w:standard_name = "ocean_s_coordinate_g1" ;
		s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
		s_w:field = "s_w, scalar" ;
	float salt(ocean_time, s_rho, eta_rho, xi_rho) ;
		salt:long_name = "salinity" ;
		salt:time = "ocean_time" ;
		salt:grid = "grid" ;
		salt:location = "face" ;
		salt:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		salt:field = "salinity, scalar, series" ;
		salt:_FillValue = 1.e+37f ;
	float sig11(ocean_time, eta_rho, xi_rho) ;
		sig11:long_name = "internal ice stress 11 component" ;
		sig11:units = "Newton meter-1" ;
		sig11:time = "ocean_time" ;
		sig11:grid = "grid" ;
		sig11:location = "face" ;
		sig11:coordinates = "lon_rho lat_rho ocean_time" ;
		sig11:field = "ice stress 11, scalar, series" ;
		sig11:_FillValue = 1.e+37f ;
	float sig12(ocean_time, eta_rho, xi_rho) ;
		sig12:long_name = "internal ice stress 12 component" ;
		sig12:units = "Newton meter-1" ;
		sig12:time = "ocean_time" ;
		sig12:grid = "grid" ;
		sig12:location = "face" ;
		sig12:coordinates = "lon_rho lat_rho ocean_time" ;
		sig12:field = "ice stress 12, scalar, series" ;
		sig12:_FillValue = 1.e+37f ;
	float sig22(ocean_time, eta_rho, xi_rho) ;
		sig22:long_name = "internal ice stress 22 component" ;
		sig22:units = "Newton meter-1" ;
		sig22:time = "ocean_time" ;
		sig22:grid = "grid" ;
		sig22:location = "face" ;
		sig22:coordinates = "lon_rho lat_rho ocean_time" ;
		sig22:field = "ice stress 22, scalar, series" ;
		sig22:_FillValue = 1.e+37f ;
	float snow_thick(ocean_time, eta_rho, xi_rho) ;
		snow_thick:long_name = "thickness of snow cover" ;
		snow_thick:units = "meter" ;
		snow_thick:time = "ocean_time" ;
		snow_thick:grid = "grid" ;
		snow_thick:location = "face" ;
		snow_thick:coordinates = "lon_rho lat_rho ocean_time" ;
		snow_thick:field = "snow thickness, scalar, series" ;
		snow_thick:_FillValue = 1.e+37f ;
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = 0, 1 ;
		spherical:flag_meanings = "Cartesian spherical" ;
	float t0mk(ocean_time, eta_rho, xi_rho) ;
		t0mk:long_name = "temperature of molecular sub-layer under ice" ;
		t0mk:units = "degrees Celsius" ;
		t0mk:time = "ocean_time" ;
		t0mk:grid = "grid" ;
		t0mk:location = "face" ;
		t0mk:coordinates = "lon_rho lat_rho ocean_time" ;
		t0mk:field = "temperature, scalar, series" ;
		t0mk:_FillValue = 1.e+37f ;
	float tau_iw(ocean_time, eta_rho, xi_rho) ;
		tau_iw:long_name = "ice-water friction velocity" ;
		tau_iw:units = "meter second-1" ;
		tau_iw:time = "ocean_time" ;
		tau_iw:grid = "grid" ;
		tau_iw:location = "face" ;
		tau_iw:coordinates = "lon_rho lat_rho ocean_time" ;
		tau_iw:field = "friction velocity, scalar, series" ;
		tau_iw:_FillValue = 1.e+37f ;
	float temp(ocean_time, s_rho, eta_rho, xi_rho) ;
		temp:long_name = "potential temperature" ;
		temp:units = "Celsius" ;
		temp:time = "ocean_time" ;
		temp:grid = "grid" ;
		temp:location = "face" ;
		temp:coordinates = "lon_rho lat_rho s_rho ocean_time" ;
		temp:field = "temperature, scalar, series" ;
		temp:_FillValue = 1.e+37f ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	float ti(ocean_time, eta_rho, xi_rho) ;
		ti:long_name = "interior ice temperature" ;
		ti:units = "degrees Celcius" ;
		ti:time = "ocean_time" ;
		ti:grid = "grid" ;
		ti:location = "face" ;
		ti:coordinates = "lon_rho lat_rho ocean_time" ;
		ti:field = "interior temperature, scalar, series" ;
		ti:_FillValue = 1.e+37f ;
	float tisrf(ocean_time, eta_rho, xi_rho) ;
		tisrf:long_name = "temperature of ice surface" ;
		tisrf:units = "degrees Celcius" ;
		tisrf:time = "ocean_time" ;
		tisrf:grid = "grid" ;
		tisrf:location = "face" ;
		tisrf:coordinates = "lon_rho lat_rho ocean_time" ;
		tisrf:field = "surface temperature, scalar, series" ;
		tisrf:_FillValue = 1.e+37f ;
	float u(ocean_time, s_rho, eta_u, xi_u) ;
		u:long_name = "u-momentum component" ;
		u:units = "meter second-1" ;
		u:time = "ocean_time" ;
		u:grid = "grid" ;
		u:location = "edge1" ;
		u:coordinates = "lon_u lat_u s_rho ocean_time" ;
		u:field = "u-velocity, scalar, series" ;
		u:_FillValue = 1.e+37f ;
	float ubar(ocean_time, eta_u, xi_u) ;
		ubar:long_name = "vertically integrated u-momentum component" ;
		ubar:units = "meter second-1" ;
		ubar:time = "ocean_time" ;
		ubar:grid = "grid" ;
		ubar:location = "edge1" ;
		ubar:coordinates = "lon_u lat_u ocean_time" ;
		ubar:field = "ubar-velocity, scalar, series" ;
		ubar:_FillValue = 1.e+37f ;
	float uice(ocean_time, eta_u, xi_u) ;
		uice:long_name = "u-component of ice velocity" ;
		uice:units = "meter second-1" ;
		uice:time = "ocean_time" ;
		uice:grid = "grid" ;
		uice:location = "edge1" ;
		uice:coordinates = "lon_u lat_u ocean_time" ;
		uice:field = "u-component of ice velocity, scalar, series" ;
		uice:_FillValue = 1.e+37f ;
	float v(ocean_time, s_rho, eta_v, xi_v) ;
		v:long_name = "v-momentum component" ;
		v:units = "meter second-1" ;
		v:time = "ocean_time" ;
		v:grid = "grid" ;
		v:location = "edge2" ;
		v:coordinates = "lon_v lat_v s_rho ocean_time" ;
		v:field = "v-velocity, scalar, series" ;
		v:_FillValue = 1.e+37f ;
	float vbar(ocean_time, eta_v, xi_v) ;
		vbar:long_name = "vertically integrated v-momentum component" ;
		vbar:units = "meter second-1" ;
		vbar:time = "ocean_time" ;
		vbar:grid = "grid" ;
		vbar:location = "edge2" ;
		vbar:coordinates = "lon_v lat_v ocean_time" ;
		vbar:field = "vbar-velocity, scalar, series" ;
		vbar:_FillValue = 1.e+37f ;
	float vice(ocean_time, eta_v, xi_v) ;
		vice:long_name = "v-component of ice velocity" ;
		vice:units = "meter second-1" ;
		vice:time = "ocean_time" ;
		vice:grid = "grid" ;
		vice:location = "edge2" ;
		vice:coordinates = "lon_v lat_v ocean_time" ;
		vice:field = "v-component of ice velocity, scalar, series" ;
		vice:_FillValue = 1.e+37f ;
	int w_L ;
		w_L:long_name = "large detritus sinking rate" ;
		w_L:units = "m d^-1" ;
	int w_S ;
		w_S:long_name = "small detritus sinking rate" ;
		w_S:units = "m d^-1" ;
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	float zeta(ocean_time, eta_rho, xi_rho) ;
		zeta:long_name = "free-surface" ;
		zeta:units = "meter" ;
		zeta:time = "ocean_time" ;
		zeta:grid = "grid" ;
		zeta:location = "face" ;
		zeta:coordinates = "lon_rho lat_rho ocean_time" ;
		zeta:field = "free-surface, scalar, series" ;
		zeta:_FillValue = 1.e+37f ;

// global attributes:
		:file = "bgcmip_banas/Out/bgcmip_banas_11_rst.nc" ;
		:format = "netCDF-3 64bit offset file" ;
		:Conventions = "CF-1.4, SGRID-0.3" ;
		:type = "ROMS/TOMS restart file" ;
		:title = "Bering Sea 10km Grid" ;
		:var_info = "../bering-Apps/Apps/Bering_BGC_variants/varinfo_banas_scaledbry.dat" ;
		:rst_file = "bgcmip_banas/Out/bgcmip_banas_11_rst.nc" ;
		:his_base = "bgcmip_banas/Out/bgcmip_banas_his" ;
		:avg_base = "bgcmip_banas/Out/bgcmip_banas_avg" ;
		:dia_base = "bgcmip_banas/Out/bgcmip_banas_dia" ;
		:sta_file = "bgcmip_banas/Out/bgcmip_banas_11_sta.nc" ;
		:grd_file = "../../ROMS_Datasets/grids/AlaskaGrids_Bering10K.nc" ;
		:ini_file = "bgcmip_banas/Out/bgcmip_banas_10_rst.nc" ;
		:tide_file = "../../ROMS_Datasets/OTPS/tides_OTPS_Bering10K.nc" ;
		:frc_file_01 = "../../ROMS_Datasets/BarrowCO2/atmo_co2_barrow_1970_2020.nc" ;
		:frc_file_02 = "../../ROMS_Datasets/Iron/ESM4_Bering10K_iron_dust_clim.nc" ;
		:frc_file_03 = "../../ROMS_Datasets/salinity/sss.clim.nc" ;
		:frc_file_04 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Pair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Pair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Pair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Pair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Pair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Pair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Pair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Pair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Pair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Pair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Pair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Pair-2020.nc" ;
		:frc_file_05 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Qair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Qair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Qair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Qair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Qair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Qair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Qair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Qair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Qair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Qair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Qair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Qair-2020.nc" ;
		:frc_file_06 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Tair-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Tair-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Tair-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Tair-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Tair-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Tair-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Tair-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Tair-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Tair-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Tair-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Tair-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Tair-2020.nc" ;
		:frc_file_07 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Uwind-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Uwind-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Uwind-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Uwind-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Uwind-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Uwind-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Uwind-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Uwind-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Uwind-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Uwind-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Uwind-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Uwind-2020.nc" ;
		:frc_file_08 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Vwind-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Vwind-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Vwind-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-Vwind-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Vwind-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Vwind-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-Vwind-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Vwind-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-Vwind-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Vwind-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-Vwind-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Vwind-2020.nc" ;
		:frc_file_09 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-rain-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-rain-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-rain-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-rain-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-rain-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-rain-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-rain-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-rain-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-rain-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-rain-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-rain-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-rain-2020.nc" ;
		:frc_file_10 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-swrad-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-swrad-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-swrad-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-swrad-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-swrad-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-swrad-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-swrad-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-swrad-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-swrad-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-swrad-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-swrad-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-swrad-2020.nc" ;
		:frc_file_11 = "../../ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-lwrad-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-lwrad-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-lwrad-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-atmos-northPacific-lwrad-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-lwrad-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-lwrad-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-lwrad-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-lwrad-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-atmos-northPacific-lwrad-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-lwrad-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-atmos-northPacific-lwrad-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-lwrad-2020.nc" ;
		:frc_file_12 = "../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2009.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2010.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2011.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2012.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2013.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2014.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2015.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2016.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2017.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2018.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2019.nc, ../../ROMS_Datasets/GloFAS/GloFAS_runoff_Bering10K_2020.nc" ;
		:frc_file_13 = "../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2009.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2010.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2011.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2012.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2013.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2014.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2015.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2016.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2017.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2018.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2019.nc, ../../ROMS_Datasets/GloFAS/GloFAS-based_nutrientflux_Bering10K_2020.nc" ;
		:bry_file_01 = "../../ROMS_Datasets/WOA2018/WOA2018_Bering10K_N30_brybgc.nc" ;
		:bry_file_02 = "../../ROMS_Datasets/CFS/2009/CFS-ocean-Bering10K-N30-bryocn-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-ocean-Bering10K-N30-bryocn-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-ocean-Bering10K-N30-bryocn-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-ocean-Bering10K-N30-bryocn-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-ocean-Bering10K-N30-bryocn-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-ocean-Bering10K-N30-bryocn-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-ocean-Bering10K-N30-bryocn-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-ocean-Bering10K-N30-bryocn-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-ocean-Bering10K-N30-bryocn-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-ocean-Bering10K-N30-bryocn-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-ocean-Bering10K-N30-bryocn-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-ocean-Bering10K-N30-bryocn-2020.nc" ;
		:bry_file_03 = "../../ROMS_Datasets/CFS/2009/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2009.nc, ../../ROMS_Datasets/CFS/2010/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2010.nc, ../../ROMS_Datasets/CFS/2011/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2011.nc, ../../ROMS_Datasets/CFS/2012/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2012.nc, ../../ROMS_Datasets/CFS/2013/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2013.nc, ../../ROMS_Datasets/CFS/2014/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2014.nc, ../../ROMS_Datasets/CFS/2015/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2015.nc, ../../ROMS_Datasets/CFS/2016/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2016.nc, ../../ROMS_Datasets/CFS/2017/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2017.nc, ../../ROMS_Datasets/CFS/2018/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2018.nc, ../../ROMS_Datasets/CFS/2019/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2019.nc, ../../ROMS_Datasets/CFS/2020/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2020.nc" ;
		:script_file = "bgcmip_banas/In/bgcmip_banas_11_ocean.in" ;
		:bpar_file = "bgcmip_banas/In/bgcmip_banas_bpar.in" ;
		:spos_file = "bgcmip_banas/In/bgcmip_banas_spos.in" ;
		:NLM_TADV = "\n",
			"ADVECTION:  HORIZONTAL   VERTICAL     \n",
			"temp:       Centered4    Centered4    \n",
			"salt:       Centered4    Centered4    \n",
			"phyto:      HSIMT        HSIMT        \n",
			"microzoo:   HSIMT        HSIMT        \n",
			"det_small:  HSIMT        HSIMT        \n",
			"det_large:  HSIMT        HSIMT        \n",
			"NH4:        HSIMT        HSIMT        \n",
			"NO3:        HSIMT        HSIMT" ;
		:NLM_LBC = "\n",
			"EDGE:        WEST   SOUTH  EAST   NORTH  \n",
			"zeta:        Che    Che    Clo    Clo    \n",
			"ubar:        Fla    Fla    Clo    Clo    \n",
			"vbar:        Fla    Fla    Clo    Clo    \n",
			"u:           RadNud RadNud Clo    Clo    \n",
			"v:           RadNud RadNud Clo    Clo    \n",
			"temp:        RadNud RadNud Clo    Clo    \n",
			"salt:        RadNud RadNud Clo    Clo    \n",
			"phyto:       RadNud RadNud Clo    Clo    \n",
			"microzoo:    RadNud RadNud Clo    Clo    \n",
			"det_small:   RadNud RadNud Clo    Clo    \n",
			"det_large:   RadNud RadNud Clo    Clo    \n",
			"NH4:         RadNud RadNud Clo    Clo    \n",
			"NO3:         RadNud RadNud Clo    Clo    \n",
			"uice:        Gra    Gra    Clo    Clo    \n",
			"vice:        Gra    Gra    Clo    Clo    \n",
			"aice:        Clo    Clo    Clo    Clo    \n",
			"hice:        Clo    Clo    Clo    Clo    \n",
			"tisrf:       Clo    Clo    Clo    Clo    \n",
			"snow_thick:  Clo    Clo    Clo    Clo    \n",
			"sig11:       Clo    Clo    Clo    Clo    \n",
			"sig12:       Clo    Clo    Clo    Clo    \n",
			"sig22:       Clo    Clo    Clo    Clo" ;
		:git_url = "git@github.com:beringnpz/roms.git" ;
		:git_rev = "cobalttweaks commit 42132fdbf454dfead62591c1ccb4f1b24400b6ab" ;
		:code_dir = "/gscratch/bumblereem/kearney/roms-kate-ice" ;
		:header_dir = "/gscratch/bumblereem/kearney/BGC_hindcasts_workdir" ;
		:header_file = "bering_10k.h" ;
		:os = "Linux" ;
		:cpu = "x86_64" ;
		:compiler_system = "ifort" ;
		:compiler_command = "/gscratch/sw/intel-201703/compilers_and_libraries_2017.2.174/linux/mpi/intel64/b" ;
		:compiler_flags = "-fp-model precise -heap-arrays -ip -O3 -traceback -check uninit -ip -O3" ;
		:tiling = "007x020" ;
		:history = "Fri Sep 22 11:02:54 2023: ncks -F -d ocean_time,2,2 /gscratch/bumblereem/kearney/BGC_hindcasts_workdir/bgcmip_banas/Out/bgcmip_banas_11_rst.nc ../ini_hindcastloop2_BIO_BANAS.nc\n",
			"ROMS/TOMS, Version 3.9, Sunday - June 25, 2023 -  7:03:52 AM" ;
		:ana_file = "ROMS/Functionals/ana_btflux.h, /gscratch/bumblereem/kearney/BGC_hindcasts_workdir/ana_psource.h, ROMS/Functionals/ana_srflux.h, ROMS/Functionals/ana_stflux.h, ROMS/Functionals/ana_aiobc.h, ROMS/Functionals/ana_hiobc.h, ROMS/Functionals/ana_hsnobc.h" ;
		:bio_file = "ROMS/Nonlinear/Biology/banas.h" ;
		:CPP_options = "BERING_10K, ADD_FSOBC, ADD_M2OBC, ALBEDO_CURVE, ANA_BPFLUX, ANA_BSFLUX, ANA_BTFLUX, ANA_PSOURCE, ANA_SPFLUX, ASSUMED_SHAPE, AVERAGES, !BOUNDARY_ALLGATHER, BULK_FLUXES, CCSM_FLUXES, COLLECT_ALLGATHER, COASTAL_ATTEN, CORE_FORCING, CURVGRID, DIAGNOSTICS_BIO, DIAGNOSTICS_TS, DIFF_GRID, DIURNAL_SRFLUX, DJ_GRADPS, DOUBLE_PRECISION, EMINUSP, ICE_ADVECT, ICE_BULK_FLUXES, ICE_EVP, ICE_MK, ICE_MODEL, ICE_MOMENTUM, ICE_SMOLAR, ICE_THERMO, LIMIT_BSTRESS, LMD_CONVEC, LMD_MIXING, LMD_NONLOCAL, LMD_RIMIX, LMD_SHAPIRO, LMD_SKPP, LONGWAVE_OUT, MASKING, MIX_GEO_TS, MIX_S_UV, MPI, NONLINEAR, NONLIN_EOS, NO_WRITE_GRID, OPTIC_MANIZZA, POT_TIDES, POWER_LAW, PROFILE, RADIATION_2D, REDUCE_ALLGATHER, RUNOFF, RST_SINGLE, SALINITY, SCORRECTION, SOLAR_SOURCE, SOLVE3D, SSH_TIDES, STATIONS, TIDES_ASTRO, TS_DIF2, UV_ADV, UV_COR, UV_U3HADVECTION, UV_SADVECTION, UV_DRAG_GRID, UV_LDRAG, UV_TIDES, UV_VIS2, UV_SMAGORINSKY, VAR_RHO_2D, VISC_GRID, VISC_3DCOEF" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
