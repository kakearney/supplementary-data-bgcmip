netcdf CFS-atmos-northPacific-Qair-1992 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:missing_value = -1.e+34 ;
		Qair:_FillValue = -1.e+34 ;
		Qair:time = "qair_time" ;
		Qair:coordinates = "lon lat" ;
		Qair:height_above_ground = 2.f ;
		Qair:long_name = "specific humidity" ;
		Qair:history = "From roms-cfs-atmos-Qair-1992" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double qair_time(qair_time) ;
		qair_time:units = "day since 1900-01-01 00:00:00" ;
		qair_time:time_origin = "01-JAN-1900 00:00:00" ;
		qair_time:axis = "T" ;
		qair_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:28:06 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1992/roms-cfs-atmos-Qair-1992.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1992/CFS-atmos-northPacific-Qair-1992.nc\n",
			"Wed Nov 20 14:00:48 2019: Time overhang added to both ends\n",
			"Wed Nov 20 14:00:40 2019: ncrcat /tmp/tp0805571f_4cc2_46eb_9c10_efd32c908067.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1992/roms-cfs-atmos-Qair-1992.nc /tmp/tpf53e9333_3a33_4a79_88de_5971ca92aacc.nc /tmp/tpa958a38b_d61f_4f29_a3e5_884644a792a9.nc\n",
			"Wed Nov 20 14:00:39 2019: ncks -F -d qair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1992/roms-cfs-atmos-Qair-1992.nc /tmp/tp0805571f_4cc2_46eb_9c10_efd32c908067.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
