netcdf CFS-atmos-northPacific-Pair-2014 {
dimensions:
	pair_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:30:46 2022: ncks -F -O -d pair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2014/roms-cfs-atmos-Pair-2014.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Pair-2014.nc\n",
			"Mon Sep 10 13:33:43 2018: Time overhang added\n",
			"Mon Sep 10 13:33:35 2018: ncrcat /tmp/tpc5839a64_b40e_49a6_8dd2_41ac94874921.nc frc/roms-cfs-atmos-Pair-2014.nc /tmp/tp9338929e_f3dc_486b_8e72_fe8a24f4c9b1.nc /tmp/tp0d3e5d33_6bf1_41ed_977c_9dae0e0fc0b5.nc\n",
			"Mon Sep 10 13:33:35 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2014.nc /tmp/tpc5839a64_b40e_49a6_8dd2_41ac94874921.nc\n",
			"Thu Sep  6 13:13:20 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2014.nc\n",
			"Thu Sep  6 13:11:15 2018: ncks -O -F -d air_time,2,1449 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2014_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2014.nc\n",
			"04-Oct-2017 18:25:09: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
