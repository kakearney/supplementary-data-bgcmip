netcdf CFS-atmos-northPacific-Vwind-1991 {
dimensions:
	wind_time = UNLIMITED ; // (1459 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:missing_value = -1.e+34 ;
		Vwind:_FillValue = -1.e+34 ;
		Vwind:time = "wind_time" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:height_above_ground1 = 10.f ;
		Vwind:long_name = "V wind" ;
		Vwind:history = "From roms-cfs-atmos-Vwind-1991" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:26:32 2022: ncks -F -O -d wind_time,2,1460 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Vwind-1991.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1991/CFS-atmos-northPacific-Vwind-1991.nc\n",
			"Wed Nov 20 13:59:17 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:59:12 2019: ncrcat /tmp/tpc7c23e2d_f92a_44ae_9dc4_787a618c64be.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Vwind-1991.nc /tmp/tp41f1ef88_8ebe_480e_a062_72f99d03aab8.nc /tmp/tpd1c68ae5_02b5_405f_9bab_8f8d342d0e21.nc\n",
			"Wed Nov 20 13:59:10 2019: ncks -F -d wind_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-Vwind-1991.nc /tmp/tpc7c23e2d_f92a_44ae_9dc4_787a618c64be.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
