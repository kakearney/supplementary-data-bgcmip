netcdf CFS-atmos-northPacific-Qair-2014 {
dimensions:
	qair_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:31:00 2022: ncks -F -O -d qair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2014/roms-cfs-atmos-Qair-2014.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-Qair-2014.nc\n",
			"Mon Sep 10 13:36:38 2018: Time overhang added\n",
			"Mon Sep 10 13:36:31 2018: ncrcat /tmp/tp30beb07e_2cc0_4179_8740_11a68fd134eb.nc frc/roms-cfs-atmos-Qair-2014.nc /tmp/tp2cf8c18a_902c_49c3_8942_901a3d1f840c.nc /tmp/tpb5fd2bfc_4641_4a58_a40b_1231373ebfb6.nc\n",
			"Mon Sep 10 13:36:30 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2014.nc /tmp/tp30beb07e_2cc0_4179_8740_11a68fd134eb.nc\n",
			"Thu Sep  6 13:23:31 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2014.nc\n",
			"Thu Sep  6 13:22:02 2018: ncks -O -F -d air_time,2,1449 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2014_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2014.nc\n",
			"04-Oct-2017 18:25:09: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
