netcdf CFS-atmos-northPacific-swrad-1996 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (366 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:43:56 2022: ncks -F -O -d srf_time,2,367 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1996/roms-cfs-atmos-swrad-1996.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1996/CFS-atmos-northPacific-swrad-1996.nc\n",
			"Mon Sep 10 14:03:42 2018: Time overhang added\n",
			"Mon Sep 10 14:03:41 2018: ncrcat /tmp/tpc355a8d5_fee0_48fc_8e7f_c0219cba2735.nc frc/roms-cfs-atmos-swrad-1996.nc /tmp/tpbc517b56_a90e_44e6_a3cf_28a4538ee307.nc /tmp/tp84ac2038_9f54_4b63_9894_fb6b5aac8e8c.nc\n",
			"Mon Sep 10 14:03:41 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-1996.nc /tmp/tpc355a8d5_fee0_48fc_8e7f_c0219cba2735.nc\n",
			"Thu Sep  6 10:01:06 2018: ncks -O -F -d srf_time,2,367 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1996_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-1996.nc\n",
			"04-Oct-2017 17:40:40: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
