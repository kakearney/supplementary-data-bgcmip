netcdf CFS-atmos-northPacific-Vwind-2011 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:05:20 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2011/roms-cfs-atmos-Vwind-2011.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-Vwind-2011.nc\n",
			"Mon Sep 10 13:45:03 2018: Time overhang added\n",
			"Mon Sep 10 13:44:55 2018: ncrcat /tmp/tp7c2f4de1_57ae_4a3a_a025_158a8057842b.nc frc/roms-cfs-atmos-Vwind-2011.nc /tmp/tpbef956c8_0549_41f5_868a_9620acc28631.nc /tmp/tp9d66ab5e_edf8_40d0_92c3_dc39d1ed5846.nc\n",
			"Mon Sep 10 13:44:54 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2011.nc /tmp/tp7c2f4de1_57ae_4a3a_a025_158a8057842b.nc\n",
			"Thu Sep  6 12:30:10 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2011_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2011.nc\n",
			"04-Oct-2017 18:15:42: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
