netcdf CFS-atmos-northPacific-Vwind-1984 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:missing_value = -1.e+34 ;
		Vwind:_FillValue = -1.e+34 ;
		Vwind:time = "wind_time" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:height_above_ground1 = 10.f ;
		Vwind:long_name = "V wind" ;
		Vwind:history = "From roms-cfs-atmos-Vwind-1984" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Thu Nov  3 15:34:58 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Vwind-1984.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1984/CFS-atmos-northPacific-Vwind-1984.nc\n",
			"Wed Nov 20 13:44:49 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:44:42 2019: ncrcat /tmp/tp4f905748_6a04_4bad_abb2_ab9b8e2f5644.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Vwind-1984.nc /tmp/tp2ef4a03a_74ce_4652_8df2_203bc320f908.nc /tmp/tp1455dcd2_fca5_43b3_bdfc_bb3a10463c4a.nc\n",
			"Wed Nov 20 13:44:40 2019: ncks -F -d wind_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Vwind-1984.nc /tmp/tp4f905748_6a04_4bad_abb2_ab9b8e2f5644.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
