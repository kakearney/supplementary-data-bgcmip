netcdf CFS-atmos-northPacific-Pair-2005 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:26 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2005/roms-cfs-atmos-Pair-2005.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2005/CFS-atmos-northPacific-Pair-2005.nc\n",
			"Mon Sep 10 13:32:33 2018: Time overhang added\n",
			"Mon Sep 10 13:32:30 2018: ncrcat /tmp/tp9135c502_e45f_4808_aa2b_0cfd27850dbd.nc frc/roms-cfs-atmos-Pair-2005.nc /tmp/tp1a28adc9_aaf4_4b4d_b972_166a0383c620.nc /tmp/tp26227935_1c5e_4345_ac03_7f7a3e6f78e8.nc\n",
			"Mon Sep 10 13:32:30 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2005.nc /tmp/tp9135c502_e45f_4808_aa2b_0cfd27850dbd.nc\n",
			"Thu Sep  6 11:17:24 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2005.nc\n",
			"Thu Sep  6 11:16:12 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2005_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2005.nc\n",
			"04-Oct-2017 18:01:29: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
