netcdf CFS-atmos-northPacific-lwrad-2015 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:46:11 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2015/roms-cfs-atmos-lwrad-2015.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2015/CFS-atmos-northPacific-lwrad-2015.nc\n",
			"Mon Sep 10 13:48:55 2018: Time overhang added\n",
			"Mon Sep 10 13:48:47 2018: ncrcat /tmp/tp8ed71f42_927b_407f_9718_84712e34bee2.nc frc/roms-cfs-atmos-lwrad-2015.nc /tmp/tpc60efb1b_1eec_4115_82eb_18d37851126f.nc /tmp/tpff38c0d5_e703_4293_a703_c97333e47f6a.nc\n",
			"Mon Sep 10 13:48:47 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2015.nc /tmp/tp8ed71f42_927b_407f_9718_84712e34bee2.nc\n",
			"Thu Sep  6 13:49:31 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2015_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2015.nc\n",
			"04-Oct-2017 18:30:21: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
