netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-2001 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:19:27 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 15:17:48 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2001/CFS-ocean-Bering10K-N30-bryocn-2001.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2001/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2001.nc\n",
			"Sat Dec 24 13:30:40 2022: ncrcat -O <>/final/2001/CFS-ocean-Bering10K-N30-bryocn-2001.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad73.nc <>/final/2001/CFS-ocean-Bering10K-N30-bryocn-2001.nc\n",
			"Wed Dec 21 13:36:24 2022: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad02.nc <>/final/2001/CFS-ocean-Bering10K-N30-bryocn-2001.nc\n",
			"Wed Dec 21 13:36:24 2022: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad01.nc\n",
			"Wed Dec 21 13:36:23 2022: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad01.nc\n",
			"Wed Dec 21 13:36:23 2022: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2001010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2001pentad01.nc\n",
			"Tue Dec 20 15:09:40 2022: CFS data added\n",
			"Tue Dec 20 15:09:11 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
