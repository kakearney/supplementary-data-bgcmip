netcdf CFS-atmos-northPacific-lwrad-2009 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:59:46 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2009/roms-cfs-atmos-lwrad-2009.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-lwrad-2009.nc\n",
			"Mon Sep 10 13:47:50 2018: Time overhang added\n",
			"Mon Sep 10 13:47:47 2018: ncrcat /tmp/tpb93d1561_fd32_47ac_bbc4_a500a928fba9.nc frc/roms-cfs-atmos-lwrad-2009.nc /tmp/tp8ab50bcf_4107_4d7c_9cf8_f3548b29dbed.nc /tmp/tp4adb8b25_7f97_41de_bf09_52b46b2cccc0.nc\n",
			"Mon Sep 10 13:47:46 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2009.nc /tmp/tpb93d1561_fd32_47ac_bbc4_a500a928fba9.nc\n",
			"Thu Sep  6 12:01:55 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2009_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2009.nc\n",
			"04-Oct-2017 18:10:10: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
