netcdf CFS-atmos-northPacific-Vwind-2020 {
dimensions:
	wind_time = UNLIMITED ; // (1448 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:missing_value = -1.e+34 ;
		Vwind:_FillValue = -1.e+34 ;
		Vwind:time = "wind_time" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:height_above_ground1 = 10.f ;
		Vwind:long_name = "V wind" ;
		Vwind:history = "From roms-cfs-atmos-Vwind-2020" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:55:46 2022: ncks -F -O -d wind_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Vwind-2020.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-Vwind-2020.nc\n",
			"Wed Jan 27 10:11:56 2021: Time overhang added to both ends\n",
			"Wed Jan 27 10:11:45 2021: ncrcat /tmp/tpe42d2e74_2506_4259_b381_fc3dacab851a.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Vwind-2020.nc /tmp/tp5714affe_7320_461f_9a2b_3c74a9d75f52.nc /tmp/tp4926c628_9c8e_4127_bd56_f28b2763b69d.nc\n",
			"Wed Jan 27 10:11:44 2021: ncks -F -d wind_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-Vwind-2020.nc /tmp/tpe42d2e74_2506_4259_b381_fc3dacab851a.nc\n",
			"FERRET V7.6  26-Jan-21" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
