netcdf CFS-atmos-northPacific-Uwind-2009 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:58:53 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2009/roms-cfs-atmos-Uwind-2009.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Uwind-2009.nc\n",
			"Mon Sep 10 13:41:42 2018: Time overhang added\n",
			"Mon Sep 10 13:41:38 2018: ncrcat /tmp/tp94958415_8952_457c_abc3_9df47cb3303e.nc frc/roms-cfs-atmos-Uwind-2009.nc /tmp/tpb574a289_2bde_4432_8d16_bc6768901de4.nc /tmp/tp7b1ee478_23f7_4b2d_8112_ad415e40f3f7.nc\n",
			"Mon Sep 10 13:41:38 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2009.nc /tmp/tp94958415_8952_457c_abc3_9df47cb3303e.nc\n",
			"Thu Sep  6 12:03:33 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2009_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2009.nc\n",
			"04-Oct-2017 18:10:30: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
