netcdf CFS-atmos-northPacific-Pair-1996 {
dimensions:
	pair_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:41:19 2022: ncks -F -O -d pair_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1996/roms-cfs-atmos-Pair-1996.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1996/CFS-atmos-northPacific-Pair-1996.nc\n",
			"Mon Sep 10 13:31:36 2018: Time overhang added\n",
			"Mon Sep 10 13:31:33 2018: ncrcat /tmp/tp5e028c6e_cfb9_4702_9fe8_8a575b8bb2a5.nc frc/roms-cfs-atmos-Pair-1996.nc /tmp/tpd1a93862_42e8_4532_971e_9fa4d183d8e5.nc /tmp/tp9b17fd89_fe40_4d6a_8b05_dc1e6cb36910.nc\n",
			"Mon Sep 10 13:31:32 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-1996.nc /tmp/tp5e028c6e_cfb9_4702_9fe8_8a575b8bb2a5.nc\n",
			"Thu Sep  6 09:56:34 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1996.nc\n",
			"Thu Sep  6 09:55:42 2018: ncks -O -F -d air_time,2,1465 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1996_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1996.nc\n",
			"04-Oct-2017 17:39:23: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
