netcdf CFS-atmos-northPacific-Uwind-2021 {
dimensions:
	wind_time = UNLIMITED ; // (1432 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:missing_value = -1.e+34 ;
		Uwind:_FillValue = -1.e+34 ;
		Uwind:time = "wind_time" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:height_above_ground1 = 10.f ;
		Uwind:long_name = "U wind" ;
		Uwind:history = "From roms-cfs-atmos-Uwind-2021" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 13:09:15 2022: ncks -F -O -d wind_time,2,1433 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2021/roms-cfs-atmos-Uwind-2021.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2021/CFS-atmos-northPacific-Uwind-2021.nc\n",
			"Fri May 06 13:51:23 2022: Time overhang added to end\n",
			"Fri May  6 13:51:15 2022: ncrcat /gscratch/bumblereem/bering10k/input/hindcast_cfs/2021/roms-cfs-atmos-Uwind-2021.nc /tmp/tp3de884e7_5983_42cf_ab5a_5fbe003a541f.nc /tmp/tp99a7f83c_e46e_43c0_bbbb_f24e6153f1e9.nc\n",
			"FERRET V7.6  20-Jan-22" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
