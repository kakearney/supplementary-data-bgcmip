netcdf CFS-atmos-northPacific-Qair-2002 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:08 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2002/roms-cfs-atmos-Qair-2002.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2002/CFS-atmos-northPacific-Qair-2002.nc\n",
			"Mon Sep 10 13:35:11 2018: Time overhang added\n",
			"Mon Sep 10 13:35:08 2018: ncrcat /tmp/tp71fb8c1b_cc74_4477_aa64_7493858f05d4.nc frc/roms-cfs-atmos-Qair-2002.nc /tmp/tpddb66103_7d1d_4465_a5ae_5a80c0b80ff7.nc /tmp/tpfec25f09_a866_461f_8cee_0733f37686c2.nc\n",
			"Mon Sep 10 13:35:07 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2002.nc /tmp/tp71fb8c1b_cc74_4477_aa64_7493858f05d4.nc\n",
			"Thu Sep  6 10:54:00 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2002.nc\n",
			"Thu Sep  6 10:52:59 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2002_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2002.nc\n",
			"04-Oct-2017 17:54:31: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
