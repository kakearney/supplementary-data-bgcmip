netcdf CFS-atmos-northPacific-Vwind-1999 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:47:48 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1999/roms-cfs-atmos-Vwind-1999.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1999/CFS-atmos-northPacific-Vwind-1999.nc\n",
			"Mon Sep 10 13:43:50 2018: Time overhang added\n",
			"Mon Sep 10 13:43:46 2018: ncrcat /tmp/tp4c16ddf3_f089_4bd3_b41a_8848185274af.nc frc/roms-cfs-atmos-Vwind-1999.nc /tmp/tp668295a6_7e3f_4f0d_9803_a5e6f74c9cd7.nc /tmp/tp161f1102_bb0f_474b_83ec_fa2962ad2a57.nc\n",
			"Mon Sep 10 13:43:46 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-1999.nc /tmp/tp4c16ddf3_f089_4bd3_b41a_8848185274af.nc\n",
			"Thu Sep  6 10:28:45 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1999_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-1999.nc\n",
			"04-Oct-2017 17:48:04: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
