netcdf CFS-atmos-northPacific-lwrad-2020 {
dimensions:
	lat = 344 ;
	lon = 588 ;
	lrf_time = UNLIMITED ; // (1447 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double lrf_time(lrf_time) ;
		lrf_time:units = "day since 1900-01-01 00:00:00" ;
		lrf_time:time_origin = "01-JAN-1900 00:00:00" ;
		lrf_time:axis = "T" ;
		lrf_time:standard_name = "time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:missing_value = -1.e+34 ;
		lwrad_down:_FillValue = -1.e+34 ;
		lwrad_down:time = "lrf_time" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:long_name = "downward longwave radiation" ;
		lwrad_down:history = "From roms-cfs-atmos-lwrad-2020" ;

// global attributes:
		:history = "Mon Oct 31 12:56:41 2022: ncks -F -O -d lrf_time,2,1448 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-lwrad-2020.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2020/CFS-atmos-northPacific-lwrad-2020.nc\n",
			"Wed Jan 27 10:12:15 2021: Time overhang added to both ends\n",
			"Wed Jan 27 10:12:05 2021: ncrcat /tmp/tpdf34d2ee_77fe_4ee9_a023_6618700071f3.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-lwrad-2020.nc /tmp/tpb10860f3_03a3_4b14_a9bd_6a505f80951e.nc /tmp/tp1834136f_d29e_45bd_892e_f1615030bd39.nc\n",
			"Wed Jan 27 10:12:04 2021: ncks -F -d lrf_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2020/roms-cfs-atmos-lwrad-2020.nc /tmp/tpdf34d2ee_77fe_4ee9_a023_6618700071f3.nc\n",
			"FERRET V7.6  26-Jan-21" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
