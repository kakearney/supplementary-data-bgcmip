netcdf CFS-atmos-northPacific-rain-1988 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double rain(rain_time, lat, lon) ;
		rain:missing_value = -1.e+34 ;
		rain:_FillValue = -1.e+34 ;
		rain:time = "rain_time" ;
		rain:coordinates = "lon lat" ;
		rain:long_name = "rainfall" ;
		rain:history = "From roms-cfs-atmos-rain-1988" ;
	double rain_time(rain_time) ;
		rain_time:units = "day since 1900-01-01 00:00:00" ;
		rain_time:time_origin = "01-JAN-1900 00:00:00" ;
		rain_time:axis = "T" ;
		rain_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:21:46 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1988/roms-cfs-atmos-rain-1988.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1988/CFS-atmos-northPacific-rain-1988.nc\n",
			"Wed Nov 20 13:53:44 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:53:37 2019: ncrcat /tmp/tpd4580fa9_571d_42b0_b4f5_cb6cd2fa2462.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1988/roms-cfs-atmos-rain-1988.nc /tmp/tp88da08ec_81ae_427e_acfd_6f78c50a5bf7.nc /tmp/tpa639c26d_5927_4a37_b69a_68f97e609d79.nc\n",
			"Wed Nov 20 13:53:35 2019: ncks -F -d rain_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1988/roms-cfs-atmos-rain-1988.nc /tmp/tpd4580fa9_571d_42b0_b4f5_cb6cd2fa2462.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
