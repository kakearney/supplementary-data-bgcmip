netcdf CFS-atmos-northPacific-swrad-2004 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (366 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:22 2022: ncks -F -O -d srf_time,2,367 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2004/roms-cfs-atmos-swrad-2004.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2004/CFS-atmos-northPacific-swrad-2004.nc\n",
			"Mon Sep 10 14:03:59 2018: Time overhang added\n",
			"Mon Sep 10 14:03:58 2018: ncrcat /tmp/tp68b79110_7830_4960_9dd5_164338f1fc14.nc frc/roms-cfs-atmos-swrad-2004.nc /tmp/tp62c84761_4566_43a4_bd55_6956cd9752b3.nc /tmp/tpc1f93205_44b1_4d24_a0e1_52df545f75d5.nc\n",
			"Mon Sep 10 14:03:58 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-2004.nc /tmp/tp68b79110_7830_4960_9dd5_164338f1fc14.nc\n",
			"Thu Sep  6 11:14:04 2018: ncks -O -F -d srf_time,2,367 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2004_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-2004.nc\n",
			"04-Oct-2017 18:00:34: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
