netcdf CFS-atmos-northPacific-Uwind-2003 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:17:09 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2003/roms-cfs-atmos-Uwind-2003.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2003/CFS-atmos-northPacific-Uwind-2003.nc\n",
			"Mon Sep 10 13:41:07 2018: Time overhang added\n",
			"Mon Sep 10 13:41:04 2018: ncrcat /tmp/tp8cfaf8a1_eb0e_4a2e_9ae6_ff798d698f13.nc frc/roms-cfs-atmos-Uwind-2003.nc /tmp/tpa02cb6f7_b84a_41c6_9edb_0b52f7d5a4f5.nc /tmp/tpd79d24e8_8b2c_4fad_b61c_127461a6b11c.nc\n",
			"Mon Sep 10 13:41:03 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2003.nc /tmp/tp8cfaf8a1_eb0e_4a2e_9ae6_ff798d698f13.nc\n",
			"Thu Sep  6 11:06:04 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2003_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2003.nc\n",
			"04-Oct-2017 17:58:25: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
