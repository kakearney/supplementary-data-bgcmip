netcdf CFS-atmos-northPacific-Qair-2010 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:00:09 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2010/roms-cfs-atmos-Qair-2010.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-Qair-2010.nc\n",
			"Mon Sep 10 13:35:54 2018: Time overhang added\n",
			"Mon Sep 10 13:35:51 2018: ncrcat /tmp/tp4303ccf6_9f77_495d_be0d_b920abd33fba.nc frc/roms-cfs-atmos-Qair-2010.nc /tmp/tpa5d0c954_fde7_4f17_9c4e_e21c3c2a3de6.nc /tmp/tp31a5ca0a_df64_4363_a710_c945a7f729cb.nc\n",
			"Mon Sep 10 13:35:51 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2010.nc /tmp/tp4303ccf6_9f77_495d_be0d_b920abd33fba.nc\n",
			"Thu Sep  6 12:08:44 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2010.nc\n",
			"Thu Sep  6 12:08:01 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2010_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2010.nc\n",
			"04-Oct-2017 18:11:27: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
