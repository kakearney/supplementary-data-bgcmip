netcdf CFS-atmos-northPacific-lwrad-2007 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:54:41 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2007/roms-cfs-atmos-lwrad-2007.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2007/CFS-atmos-northPacific-lwrad-2007.nc\n",
			"Mon Sep 10 13:47:39 2018: Time overhang added\n",
			"Mon Sep 10 13:47:35 2018: ncrcat /tmp/tp9abe9efc_050c_4da7_b6b8_48cbc3113fd1.nc frc/roms-cfs-atmos-lwrad-2007.nc /tmp/tp577795cd_15bf_4a02_aad2_9ca613d1d982.nc /tmp/tpb48d3011_77ba_42a4_8ca9_27537ae2527a.nc\n",
			"Mon Sep 10 13:47:35 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2007.nc /tmp/tp9abe9efc_050c_4da7_b6b8_48cbc3113fd1.nc\n",
			"Thu Sep  6 11:45:24 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2007_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2007.nc\n",
			"04-Oct-2017 18:06:10: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
