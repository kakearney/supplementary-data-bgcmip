netcdf CFS-atmos-northPacific-rain-1998 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:46:41 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1998/roms-cfs-atmos-rain-1998.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1998/CFS-atmos-northPacific-rain-1998.nc\n",
			"Mon Sep 10 13:50:01 2018: Time overhang added\n",
			"Mon Sep 10 13:49:57 2018: ncrcat /tmp/tp3520cbea_0843_4c7b_b55f_3d583357c1c2.nc frc/roms-cfs-atmos-rain-1998.nc /tmp/tp9c3ed9f3_08ee_4981_a4f9_604b7001dff6.nc /tmp/tpb5fbc8f1_baa5_4e9a_968a_3e3cf7b1954c.nc\n",
			"Mon Sep 10 13:49:56 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-1998.nc /tmp/tp3520cbea_0843_4c7b_b55f_3d583357c1c2.nc\n",
			"Thu Sep  6 10:17:31 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1998_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-1998.nc\n",
			"04-Oct-2017 17:46:18: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
