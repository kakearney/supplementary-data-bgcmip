netcdf CFS-atmos-northPacific-Tair-2005 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:39 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2005/roms-cfs-atmos-Tair-2005.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2005/CFS-atmos-northPacific-Tair-2005.nc\n",
			"Mon Sep 10 13:38:23 2018: Time overhang added\n",
			"Mon Sep 10 13:38:19 2018: ncrcat /tmp/tp23298660_ab37_4a99_85a0_c27a835ae52c.nc frc/roms-cfs-atmos-Tair-2005.nc /tmp/tped03360a_c147_41bf_b5e2_bfd3c82b46ec.nc /tmp/tp015a2204_64d3_4288_9dbf_b21a33f918ee.nc\n",
			"Mon Sep 10 13:38:19 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2005.nc /tmp/tp23298660_ab37_4a99_85a0_c27a835ae52c.nc\n",
			"Thu Sep  6 11:19:13 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2005.nc\n",
			"Thu Sep  6 11:18:04 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2005_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2005.nc\n",
			"04-Oct-2017 18:01:29: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
