netcdf CFS-atmos-northPacific-Uwind-2005 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:46 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2005/roms-cfs-atmos-Uwind-2005.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2005/CFS-atmos-northPacific-Uwind-2005.nc\n",
			"Mon Sep 10 13:41:18 2018: Time overhang added\n",
			"Mon Sep 10 13:41:15 2018: ncrcat /tmp/tpda7d79fe_ed01_4d14_8a0d_dd9a9e8d939e.nc frc/roms-cfs-atmos-Uwind-2005.nc /tmp/tpe880b5a4_6221_42d3_a743_cbf14c493524.nc /tmp/tp65f8293b_783e_4b19_87ab_9a2c8862c336.nc\n",
			"Mon Sep 10 13:41:14 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2005.nc /tmp/tpda7d79fe_ed01_4d14_8a0d_dd9a9e8d939e.nc\n",
			"Thu Sep  6 11:23:51 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2005_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2005.nc\n",
			"04-Oct-2017 18:02:37: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
