netcdf CFS-atmos-northPacific-Tair-2009 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:58:14 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2009/roms-cfs-atmos-Tair-2009.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2009/CFS-atmos-northPacific-Tair-2009.nc\n",
			"Mon Sep 10 13:38:45 2018: Time overhang added\n",
			"Mon Sep 10 13:38:41 2018: ncrcat /tmp/tpd78918a4_ff51_4fb5_9959_8c2630562a06.nc frc/roms-cfs-atmos-Tair-2009.nc /tmp/tpfa0a8a7b_32f8_407e_ab8f_5e5e74908153.nc /tmp/tp96cd0ba7_91fc_417e_8f9c_95c8b55ae201.nc\n",
			"Mon Sep 10 13:38:41 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2009.nc /tmp/tpd78918a4_ff51_4fb5_9959_8c2630562a06.nc\n",
			"Thu Sep  6 11:59:52 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2009.nc\n",
			"Thu Sep  6 11:59:00 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2009_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2009.nc\n",
			"04-Oct-2017 18:09:27: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
