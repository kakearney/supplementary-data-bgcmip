netcdf CFS-atmos-northPacific-lwrad-2005 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:52:01 2022: ncks -F -O -d lrf_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2005/roms-cfs-atmos-lwrad-2005.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2005/CFS-atmos-northPacific-lwrad-2005.nc\n",
			"Mon Sep 10 13:47:28 2018: Time overhang added\n",
			"Mon Sep 10 13:47:24 2018: ncrcat /tmp/tp2f00758c_23f6_4042_835b_5e8741be0b8d.nc frc/roms-cfs-atmos-lwrad-2005.nc /tmp/tp1c9af75a_419d_4494_ba7e_55cf518f7ea0.nc /tmp/tpccf2ac22_4a99_482c_a442_c60ab3e26ad8.nc\n",
			"Mon Sep 10 13:47:24 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2005.nc /tmp/tp2f00758c_23f6_4042_835b_5e8741be0b8d.nc\n",
			"Thu Sep  6 11:21:38 2018: ncks -O -F -d lrf_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2005_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2005.nc\n",
			"04-Oct-2017 18:02:15: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
