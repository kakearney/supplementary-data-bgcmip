netcdf CFS-atmos-northPacific-lwrad-2000 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	lrf_time = UNLIMITED ; // (1464 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:49:18 2022: ncks -F -O -d lrf_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2000/roms-cfs-atmos-lwrad-2000.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2000/CFS-atmos-northPacific-lwrad-2000.nc\n",
			"Mon Sep 10 13:46:59 2018: Time overhang added\n",
			"Mon Sep 10 13:46:56 2018: ncrcat /tmp/tp21e208e1_93d0_4cc4_81fa_0affcde6332e.nc frc/roms-cfs-atmos-lwrad-2000.nc /tmp/tpd18f0fae_b9fc_4021_bc27_22900971b6cc.nc /tmp/tp85f44114_52da_4174_b533_0825f8af7b0f.nc\n",
			"Mon Sep 10 13:46:55 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2000.nc /tmp/tp21e208e1_93d0_4cc4_81fa_0affcde6332e.nc\n",
			"Thu Sep  6 10:34:58 2018: ncks -O -F -d lrf_time,2,1465 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2000_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2000.nc\n",
			"04-Oct-2017 17:50:05: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
