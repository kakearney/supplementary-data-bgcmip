netcdf CFS-atmos-northPacific-Pair-1999 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:46:51 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1999/roms-cfs-atmos-Pair-1999.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1999/CFS-atmos-northPacific-Pair-1999.nc\n",
			"Mon Sep 10 13:32:00 2018: Time overhang added\n",
			"Mon Sep 10 13:31:57 2018: ncrcat /tmp/tp7607fba1_4308_4666_9101_fa44f3d6fd23.nc frc/roms-cfs-atmos-Pair-1999.nc /tmp/tpf46e07b7_fc43_44b7_8bae_225bfbf5463d.nc /tmp/tpc18d468e_bddc_424a_8ddc_f640c4027e0e.nc\n",
			"Mon Sep 10 13:31:57 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-1999.nc /tmp/tp7607fba1_4308_4666_9101_fa44f3d6fd23.nc\n",
			"Thu Sep  6 10:21:16 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1999.nc\n",
			"Thu Sep  6 10:20:07 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1999_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1999.nc\n",
			"04-Oct-2017 17:46:41: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
