netcdf CFS-atmos-northPacific-lwrad-2014 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	lrf_time = UNLIMITED ; // (1448 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double lrf_time(lrf_time) ;
		lrf_time:long_name = "forcing time" ;
		lrf_time:units = "days since 1900-01-01 00:00:00" ;
		lrf_time:time = "lrf_time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:long_name = "downwelling longwave radiation flux" ;
		lwrad_down:units = "watt meter-2" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:time = "lrf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:33:48 2022: ncks -F -O -d lrf_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2014/roms-cfs-atmos-lwrad-2014.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2014/CFS-atmos-northPacific-lwrad-2014.nc\n",
			"Mon Sep 10 13:48:43 2018: Time overhang added\n",
			"Mon Sep 10 13:48:35 2018: ncrcat /tmp/tpec65d11f_c058_4c5c_aac8_843e21c443a1.nc frc/roms-cfs-atmos-lwrad-2014.nc /tmp/tp4e017053_beee_4669_9434_f3a1f459cb59.nc /tmp/tp43767a85_52f8_416d_bd7e_8925fdb26b3e.nc\n",
			"Mon Sep 10 13:48:34 2018: ncks -F -d lrf_time,1,1 frc/roms-cfs-atmos-lwrad-2014.nc /tmp/tpec65d11f_c058_4c5c_aac8_843e21c443a1.nc\n",
			"Thu Sep  6 13:26:36 2018: ncks -O -F -d lrf_time,2,1449 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2014_lwrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-lwrad-2014.nc\n",
			"04-Oct-2017 18:26:37: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
