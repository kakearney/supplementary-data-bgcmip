netcdf CFS-atmos-northPacific-lwrad-2018 {
dimensions:
	lat = 344 ;
	lon = 588 ;
	lrf_time = UNLIMITED ; // (1452 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double lrf_time(lrf_time) ;
		lrf_time:units = "day since 1900-01-01 00:00:00" ;
		lrf_time:time_origin = "01-JAN-1900 00:00:00" ;
		lrf_time:axis = "T" ;
		lrf_time:standard_name = "time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:missing_value = -1.e+34 ;
		lwrad_down:_FillValue = -1.e+34 ;
		lwrad_down:time = "lrf_time" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:long_name = "downward longwave radiation" ;
		lwrad_down:history = "From roms-cfs-atmos-lwrad-2018" ;

// global attributes:
		:history = "Mon Oct 31 12:26:10 2022: ncks -F -O -d lrf_time,2,1453 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-lwrad-2018.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-lwrad-2018.nc\n",
			"Thu May 30 20:49:42 2019: Time overhang added\n",
			"Thu May 30 20:49:35 2019: ncrcat /tmp/tp0adc19db_eeb7_4d28_b52a_1d4accf3f2ec.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-lwrad-2018.nc /tmp/tpa7e78796_3db4_4285_a170_eb65975ccc0a.nc /tmp/tp85467358_c7a1_4e17_86a4_fd463686702e.nc\n",
			"Thu May 30 20:49:35 2019: ncks -F -d lrf_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-lwrad-2018.nc /tmp/tp0adc19db_eeb7_4d28_b52a_1d4accf3f2ec.nc\n",
			"FERRET V7.4  29-May-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
