netcdf CFS-atmos-northPacific-Qair-1998 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:44:56 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1998/roms-cfs-atmos-Qair-1998.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1998/CFS-atmos-northPacific-Qair-1998.nc\n",
			"Mon Sep 10 13:34:49 2018: Time overhang added\n",
			"Mon Sep 10 13:34:45 2018: ncrcat /tmp/tp673d54bf_3248_4ff7_b92d_742a1b218f18.nc frc/roms-cfs-atmos-Qair-1998.nc /tmp/tp4b4f9c58_ca2a_4a9d_8704_0607a39c9f8b.nc /tmp/tpe16df62d_2a6e_46c1_b96e_c385a9825bd9.nc\n",
			"Mon Sep 10 13:34:45 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-1998.nc /tmp/tp673d54bf_3248_4ff7_b92d_742a1b218f18.nc\n",
			"Thu Sep  6 10:16:20 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-1998.nc\n",
			"Thu Sep  6 10:15:37 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1998_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-1998.nc\n",
			"04-Oct-2017 17:44:14: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
