netcdf CFS-atmos-northPacific-Pair-2004 {
dimensions:
	pair_time = UNLIMITED ; // (1464 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:50:35 2022: ncks -F -O -d pair_time,2,1465 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2004/roms-cfs-atmos-Pair-2004.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2004/CFS-atmos-northPacific-Pair-2004.nc\n",
			"Mon Sep 10 13:32:28 2018: Time overhang added\n",
			"Mon Sep 10 13:32:25 2018: ncrcat /tmp/tpc4560279_6cf1_40a2_b815_2f608aec0735.nc frc/roms-cfs-atmos-Pair-2004.nc /tmp/tp1dc9add2_02e2_45fb_a43f_43cd8092a613.nc /tmp/tp9f2d8c2e_a96c_4788_a91f_f9d3cc8e4ca7.nc\n",
			"Mon Sep 10 13:32:25 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2004.nc /tmp/tpc4560279_6cf1_40a2_b815_2f608aec0735.nc\n",
			"Thu Sep  6 11:08:47 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2004.nc\n",
			"Thu Sep  6 11:07:50 2018: ncks -O -F -d air_time,2,1465 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2004_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2004.nc\n",
			"04-Oct-2017 17:59:35: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
