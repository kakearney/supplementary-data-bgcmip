netcdf CFS-atmos-northPacific-Qair-2001 {
dimensions:
	qair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Qair(qair_time, lat, lon) ;
		Qair:long_name = "surface air relative humidity" ;
		Qair:units = "kg/kg" ;
		Qair:coordinates = "lon lat" ;
		Qair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double qair_time(qair_time) ;
		qair_time:long_name = "forcing time" ;
		qair_time:units = "days since 1900-01-01 00:00:00" ;
		qair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:49:39 2022: ncks -F -O -d qair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2001/roms-cfs-atmos-Qair-2001.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2001/CFS-atmos-northPacific-Qair-2001.nc\n",
			"Mon Sep 10 13:35:06 2018: Time overhang added\n",
			"Mon Sep 10 13:35:02 2018: ncrcat /tmp/tp81e11c91_fd1c_4859_96be_b518c1e78ba6.nc frc/roms-cfs-atmos-Qair-2001.nc /tmp/tp5cb112fa_cc65_4f2e_8908_8a90f0a61c08.nc /tmp/tpf07685e4_fdb6_405e_b21a_7377d412ec78.nc\n",
			"Mon Sep 10 13:35:02 2018: ncks -F -d qair_time,1,1 frc/roms-cfs-atmos-Qair-2001.nc /tmp/tp81e11c91_fd1c_4859_96be_b518c1e78ba6.nc\n",
			"Thu Sep  6 10:43:37 2018: ncrename -d air_time,qair_time -v air_time,qair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2001.nc\n",
			"Thu Sep  6 10:42:39 2018: ncks -O -F -d air_time,2,1461 -v Qair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2001_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Qair-2001.nc\n",
			"04-Oct-2017 17:51:47: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
