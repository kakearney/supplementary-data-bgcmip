netcdf CFS-atmos-northPacific-Uwind-1986 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:missing_value = -1.e+34 ;
		Uwind:_FillValue = -1.e+34 ;
		Uwind:time = "wind_time" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:height_above_ground1 = 10.f ;
		Uwind:long_name = "U wind" ;
		Uwind:history = "From roms-cfs-atmos-Uwind-1986" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double wind_time(wind_time) ;
		wind_time:units = "day since 1900-01-01 00:00:00" ;
		wind_time:time_origin = "01-JAN-1900 00:00:00" ;
		wind_time:axis = "T" ;
		wind_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:19:44 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-Uwind-1986.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1986/CFS-atmos-northPacific-Uwind-1986.nc\n",
			"Wed Nov 20 13:48:33 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:48:26 2019: ncrcat /tmp/tp894cb699_511c_404e_a9a2_0abbdf49b86f.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-Uwind-1986.nc /tmp/tpe2ee7fc9_cd56_4338_9147_394fa08c8c4f.nc /tmp/tp7177e4de_448b_4927_9784_44708664650b.nc\n",
			"Wed Nov 20 13:48:24 2019: ncks -F -d wind_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1986/roms-cfs-atmos-Uwind-1986.nc /tmp/tp894cb699_511c_404e_a9a2_0abbdf49b86f.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
