netcdf CFS-atmos-northPacific-swrad-2010 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	srf_time = UNLIMITED ; // (365 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double srf_time(srf_time) ;
		srf_time:long_name = "forcing time" ;
		srf_time:units = "days since 1900-01-01 00:00:00" ;
		srf_time:time = "srf_time" ;
	double swrad(srf_time, lat, lon) ;
		swrad:long_name = "solar shortwave radiation flux" ;
		swrad:units = "watt meter-2" ;
		swrad:coordinates = "lon lat" ;
		swrad:time = "srf_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:02:16 2022: ncks -F -O -d srf_time,2,366 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2010/roms-cfs-atmos-swrad-2010.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2010/CFS-atmos-northPacific-swrad-2010.nc\n",
			"Mon Sep 10 14:04:13 2018: Time overhang added\n",
			"Mon Sep 10 14:04:12 2018: ncrcat /tmp/tp7a2b5d81_efbe_4898_8536_3509053020c0.nc frc/roms-cfs-atmos-swrad-2010.nc /tmp/tp1e6e315d_d391_4bab_900f_d090d963a2c1.nc /tmp/tp00e67687_c0b5_40cf_bb7e_9345679354db.nc\n",
			"Mon Sep 10 14:04:11 2018: ncks -F -d srf_time,1,1 frc/roms-cfs-atmos-swrad-2010.nc /tmp/tp7a2b5d81_efbe_4898_8536_3509053020c0.nc\n",
			"Thu Sep  6 12:10:38 2018: ncks -O -F -d srf_time,2,366 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2010_swrad.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-swrad-2010.nc\n",
			"04-Oct-2017 18:12:26: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
