netcdf CFS-atmos-northPacific-rain-2006 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:53:07 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2006/roms-cfs-atmos-rain-2006.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2006/CFS-atmos-northPacific-rain-2006.nc\n",
			"Mon Sep 10 13:50:53 2018: Time overhang added\n",
			"Mon Sep 10 13:50:49 2018: ncrcat /tmp/tpa5ee6675_0791_4abf_b4b5_134b673cb41c.nc frc/roms-cfs-atmos-rain-2006.nc /tmp/tpe847526d_ceb5_4854_93db_329f75999010.nc /tmp/tp0907a7fd_8b20_4857_a1ac_b36c8bd08031.nc\n",
			"Mon Sep 10 13:50:49 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2006.nc /tmp/tpa5ee6675_0791_4abf_b4b5_134b673cb41c.nc\n",
			"Thu Sep  6 11:35:05 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2006_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2006.nc\n",
			"04-Oct-2017 18:05:09: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
