netcdf CFS-atmos-northPacific-Uwind-2002 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Uwind(wind_time, lat, lon) ;
		Uwind:long_name = "surface u-wind component" ;
		Uwind:units = "meter second-1" ;
		Uwind:coordinates = "lon lat" ;
		Uwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:22 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2002/roms-cfs-atmos-Uwind-2002.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2002/CFS-atmos-northPacific-Uwind-2002.nc\n",
			"Mon Sep 10 13:41:02 2018: Time overhang added\n",
			"Mon Sep 10 13:40:58 2018: ncrcat /tmp/tpb99aea9e_b3d1_4143_8f96_38af0360a9b3.nc frc/roms-cfs-atmos-Uwind-2002.nc /tmp/tp8aa9d998_e24c_4a42_9772_fecac400a3cd.nc /tmp/tpa7a5df7f_d51a_4896_8060_e1de75515470.nc\n",
			"Mon Sep 10 13:40:58 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Uwind-2002.nc /tmp/tpb99aea9e_b3d1_4143_8f96_38af0360a9b3.nc\n",
			"Thu Sep  6 10:56:58 2018: ncks -O -F -d wind_time,2,1461 -v Uwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2002_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Uwind-2002.nc\n",
			"04-Oct-2017 17:56:02: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
