netcdf WOA2018_Bering10K_N30_brybgc.padded {
dimensions:
	bio_time = UNLIMITED ; // (14 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double Fe_east(bio_time, s_rho, eta_rho) ;
		Fe_east:long_name = "dissolved iron, eastern boundary condition" ;
		Fe_east:unit = "nmol/L" ;
		Fe_east:time = "bio_time" ;
		Fe_east:_FillValue = 1.e+36 ;
		Fe_east:cell_methods = "bio_time: mean" ;
	double Fe_south(bio_time, s_rho, xi_rho) ;
		Fe_south:long_name = "dissolved iron, southern boundary condition" ;
		Fe_south:unit = "nmol/L" ;
		Fe_south:time = "bio_time" ;
		Fe_south:_FillValue = 1.e+36 ;
		Fe_south:cell_methods = "bio_time: mean" ;
	double Fe_west(bio_time, s_rho, eta_rho) ;
		Fe_west:long_name = "dissolved iron, western boundary condition" ;
		Fe_west:unit = "nmol/L" ;
		Fe_west:time = "bio_time" ;
		Fe_west:_FillValue = 1.e+36 ;
		Fe_west:cell_methods = "bio_time: mean" ;
	double NH4_east(bio_time, s_rho, eta_rho) ;
		NH4_east:long_name = "ammonium, eastern boundary condition" ;
		NH4_east:unit = "umol/kg" ;
		NH4_east:time = "bio_time" ;
		NH4_east:_FillValue = 1.e+36 ;
		NH4_east:cell_methods = "bio_time: mean" ;
	double NH4_south(bio_time, s_rho, xi_rho) ;
		NH4_south:long_name = "ammonium, southern boundary condition" ;
		NH4_south:unit = "umol/kg" ;
		NH4_south:time = "bio_time" ;
		NH4_south:_FillValue = 1.e+36 ;
		NH4_south:cell_methods = "bio_time: mean" ;
	double NH4_west(bio_time, s_rho, eta_rho) ;
		NH4_west:long_name = "ammonium, western boundary condition" ;
		NH4_west:unit = "umol/kg" ;
		NH4_west:time = "bio_time" ;
		NH4_west:_FillValue = 1.e+36 ;
		NH4_west:cell_methods = "bio_time: mean" ;
	double NO3_east(bio_time, s_rho, eta_rho) ;
		NO3_east:long_name = "nitrate, eastern boundary condition" ;
		NO3_east:unit = "umol/kg" ;
		NO3_east:time = "bio_time" ;
		NO3_east:_FillValue = 1.e+36 ;
		NO3_east:cell_methods = "bio_time: mean" ;
	double NO3_south(bio_time, s_rho, xi_rho) ;
		NO3_south:long_name = "nitrate, southern boundary condition" ;
		NO3_south:unit = "umol/kg" ;
		NO3_south:time = "bio_time" ;
		NO3_south:_FillValue = 1.e+36 ;
		NO3_south:cell_methods = "bio_time: mean" ;
	double NO3_west(bio_time, s_rho, eta_rho) ;
		NO3_west:long_name = "nitrate, western boundary condition" ;
		NO3_west:unit = "umol/kg" ;
		NO3_west:time = "bio_time" ;
		NO3_west:_FillValue = 1.e+36 ;
		NO3_west:cell_methods = "bio_time: mean" ;
	double PO4_east(bio_time, s_rho, eta_rho) ;
		PO4_east:long_name = "phosphate, eastern boundary condition" ;
		PO4_east:unit = "umol/kg" ;
		PO4_east:time = "bio_time" ;
		PO4_east:_FillValue = 1.e+36 ;
		PO4_east:cell_methods = "bio_time: mean" ;
	double PO4_south(bio_time, s_rho, xi_rho) ;
		PO4_south:long_name = "phosphate, southern boundary condition" ;
		PO4_south:unit = "umol/kg" ;
		PO4_south:time = "bio_time" ;
		PO4_south:_FillValue = 1.e+36 ;
		PO4_south:cell_methods = "bio_time: mean" ;
	double PO4_west(bio_time, s_rho, eta_rho) ;
		PO4_west:long_name = "phosphate, western boundary condition" ;
		PO4_west:unit = "umol/kg" ;
		PO4_west:time = "bio_time" ;
		PO4_west:_FillValue = 1.e+36 ;
		PO4_west:cell_methods = "bio_time: mean" ;
	double SiO4_east(bio_time, s_rho, eta_rho) ;
		SiO4_east:long_name = "silicate, eastern boundary condition" ;
		SiO4_east:unit = "umol/kg" ;
		SiO4_east:time = "bio_time" ;
		SiO4_east:_FillValue = 1.e+36 ;
		SiO4_east:cell_methods = "bio_time: mean" ;
	double SiO4_south(bio_time, s_rho, xi_rho) ;
		SiO4_south:long_name = "silicate, southern boundary condition" ;
		SiO4_south:unit = "umol/kg" ;
		SiO4_south:time = "bio_time" ;
		SiO4_south:_FillValue = 1.e+36 ;
		SiO4_south:cell_methods = "bio_time: mean" ;
	double SiO4_west(bio_time, s_rho, eta_rho) ;
		SiO4_west:long_name = "silicate, western boundary condition" ;
		SiO4_west:unit = "umol/kg" ;
		SiO4_west:time = "bio_time" ;
		SiO4_west:_FillValue = 1.e+36 ;
		SiO4_west:cell_methods = "bio_time: mean" ;
	double bio_time(bio_time) ;
		bio_time:long_name = "time, climatological" ;
		bio_time:units = "days" ;
		bio_time:cycle_length = 365.25 ;
		bio_time:cell_methods = "bio_time: mean" ;
	double ones_east(bio_time, s_rho, eta_rho) ;
		ones_east:long_name = "generic tracer, eastern boundary condition" ;
		ones_east:unit = "tracer units" ;
		ones_east:time = "bio_time" ;
		ones_east:_FillValue = 1.e+36 ;
		ones_east:cell_methods = "bio_time: mean" ;
	double ones_south(bio_time, s_rho, xi_rho) ;
		ones_south:long_name = "generic tracer, southern boundary condition" ;
		ones_south:unit = "tracer units" ;
		ones_south:time = "bio_time" ;
		ones_south:_FillValue = 1.e+36 ;
		ones_south:cell_methods = "bio_time: mean" ;
	double ones_west(bio_time, s_rho, eta_rho) ;
		ones_west:long_name = "generic tracer, western boundary condition" ;
		ones_west:unit = "tracer units" ;
		ones_west:time = "bio_time" ;
		ones_west:_FillValue = 1.e+36 ;
		ones_west:cell_methods = "bio_time: mean" ;
	double oxygen_east(bio_time, s_rho, eta_rho) ;
		oxygen_east:long_name = "oxygen, eastern boundary condition" ;
		oxygen_east:unit = "umol/kg" ;
		oxygen_east:time = "bio_time" ;
		oxygen_east:_FillValue = 1.e+36 ;
		oxygen_east:cell_methods = "bio_time: mean" ;
	double oxygen_south(bio_time, s_rho, xi_rho) ;
		oxygen_south:long_name = "oxygen, southern boundary condition" ;
		oxygen_south:unit = "umol/kg" ;
		oxygen_south:time = "bio_time" ;
		oxygen_south:_FillValue = 1.e+36 ;
		oxygen_south:cell_methods = "bio_time: mean" ;
	double oxygen_west(bio_time, s_rho, eta_rho) ;
		oxygen_west:long_name = "oxygen, western boundary condition" ;
		oxygen_west:unit = "umol/kg" ;
		oxygen_west:time = "bio_time" ;
		oxygen_west:_FillValue = 1.e+36 ;
		oxygen_west:cell_methods = "bio_time: mean" ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Mon Mar 13 14:14:45 2023: Interpolated values to cycle_length time break to prevent ROMS restart issues\n",
			"Mon Mar 13 14:14:40 2023: ncrcat -O WOA2018_Bering10K_N30_brybgc_edgeinterp1.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/WOA2018/WOA2018_Bering10K_N30_brybgc.nc WOA2018_Bering10K_N30_brybgc_edgeinterp2.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/WOA2018/WOA2018_Bering10K_N30_brybgc.nc\n",
			"Mon Mar 13 14:14:39 2023: ncks -F -d bio_time,1,1 /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/WOA2018/WOA2018_Bering10K_N30_brybgc.nc WOA2018_Bering10K_N30_brybgc_edgeinterp1.nc\n",
			"Wed Jan 25 11:49:29 2023: BGC data added: NO3, PO4, O2, SiO4: World Ocean Atlas 2018 objective analysis mean (monthly surface, annual deep); Fe: Huang et al., 2022 climatology + GOANPZ analytical\n",
			"Wed Jan 25 11:49:25 2023: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
