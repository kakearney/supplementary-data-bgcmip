netcdf CFS-atmos-northPacific-Tair-2001 {
dimensions:
	tair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:49:46 2022: ncks -F -O -d tair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2001/roms-cfs-atmos-Tair-2001.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2001/CFS-atmos-northPacific-Tair-2001.nc\n",
			"Mon Sep 10 13:38:01 2018: Time overhang added\n",
			"Mon Sep 10 13:37:58 2018: ncrcat /tmp/tpc4245685_8012_4c01_8284_c4e378827ef0.nc frc/roms-cfs-atmos-Tair-2001.nc /tmp/tpe1f66910_0298_4c04_b161_9df230ff74d0.nc /tmp/tp05868eeb_7bf0_4e7c_9103_4b48c04cad70.nc\n",
			"Mon Sep 10 13:37:57 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2001.nc /tmp/tpc4245685_8012_4c01_8284_c4e378827ef0.nc\n",
			"Thu Sep  6 10:42:04 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2001.nc\n",
			"Thu Sep  6 10:40:51 2018: ncks -O -F -d air_time,2,1461 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2001_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2001.nc\n",
			"04-Oct-2017 17:51:47: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
