netcdf CFS-atmos-northPacific-lwrad-1991 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	lrf_time = UNLIMITED ; // (1459 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double lrf_time(lrf_time) ;
		lrf_time:units = "day since 1900-01-01 00:00:00" ;
		lrf_time:time_origin = "01-JAN-1900 00:00:00" ;
		lrf_time:axis = "T" ;
		lrf_time:standard_name = "time" ;
	double lwrad_down(lrf_time, lat, lon) ;
		lwrad_down:missing_value = -1.e+34 ;
		lwrad_down:_FillValue = -1.e+34 ;
		lwrad_down:time = "lrf_time" ;
		lwrad_down:coordinates = "lon lat" ;
		lwrad_down:long_name = "downward longwave radiation" ;
		lwrad_down:history = "From roms-cfs-atmos-lwrad-1991" ;

// global attributes:
		:history = "Fri Oct 28 16:27:21 2022: ncks -F -O -d lrf_time,2,1460 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-lwrad-1991.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1991/CFS-atmos-northPacific-lwrad-1991.nc\n",
			"Wed Nov 20 13:59:29 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:59:24 2019: ncrcat /tmp/tp456ea9cb_b4d3_4807_99a7_d01298c892bf.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-lwrad-1991.nc /tmp/tpeb2c3bbb_e855_49db_b068_40b61cc8ff7b.nc /tmp/tpbb660900_707c_493a_b57f_ad4e674ec665.nc\n",
			"Wed Nov 20 13:59:22 2019: ncks -F -d lrf_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1991/roms-cfs-atmos-lwrad-1991.nc /tmp/tp456ea9cb_b4d3_4807_99a7_d01298c892bf.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
