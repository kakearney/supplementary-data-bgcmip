netcdf CFS-atmos-northPacific-rain-2001 {
dimensions:
	lat = 224 ;
	lon = 384 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:50:24 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2001/roms-cfs-atmos-rain-2001.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2001/CFS-atmos-northPacific-rain-2001.nc\n",
			"Mon Sep 10 13:50:18 2018: Time overhang added\n",
			"Mon Sep 10 13:50:14 2018: ncrcat /tmp/tpb307e1bf_7c4d_47a9_bb62_3a027c2402bf.nc frc/roms-cfs-atmos-rain-2001.nc /tmp/tp35bc8396_5bf9_472f_94a5_2bdfaabf743e.nc /tmp/tp10a3f684_7a64_4656_b429_ea689b9fc72e.nc\n",
			"Mon Sep 10 13:50:14 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2001.nc /tmp/tpb307e1bf_7c4d_47a9_bb62_3a027c2402bf.nc\n",
			"Thu Sep  6 10:45:18 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2001_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2001.nc\n",
			"04-Oct-2017 17:54:07: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
