netcdf CFS-atmos-northPacific-Tair-2016 {
dimensions:
	tair_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Tair(tair_time, lat, lon) ;
		Tair:long_name = "surface air temperature" ;
		Tair:units = "Celsius" ;
		Tair:coordinates = "lon lat" ;
		Tair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double tair_time(tair_time) ;
		tair_time:long_name = "forcing time" ;
		tair_time:units = "days since 1900-01-01 00:00:00" ;
		tair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Mon Oct 31 11:55:00 2022: ncks -F -O -d tair_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2016/roms-cfs-atmos-Tair-2016.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2016/CFS-atmos-northPacific-Tair-2016.nc\n",
			"Mon Sep 10 13:39:56 2018: Time overhang added\n",
			"Mon Sep 10 13:39:49 2018: ncrcat /tmp/tp147ec2b5_cb76_4e83_8922_c41cc4cc7b22.nc frc/roms-cfs-atmos-Tair-2016.nc /tmp/tpbf5e9b24_e294_4f62_af6f_e0675df07226.nc /tmp/tpc55bfda5_318f_491c_9d16_f6997e0775e2.nc\n",
			"Mon Sep 10 13:39:48 2018: ncks -F -d tair_time,1,1 frc/roms-cfs-atmos-Tair-2016.nc /tmp/tp147ec2b5_cb76_4e83_8922_c41cc4cc7b22.nc\n",
			"Thu Sep  6 14:05:42 2018: ncrename -d air_time,tair_time -v air_time,tair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2016.nc\n",
			"Thu Sep  6 14:03:21 2018: ncks -O -F -d air_time,2,1449 -v Tair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2016_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Tair-2016.nc\n",
			"04-Oct-2017 18:32:42: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
