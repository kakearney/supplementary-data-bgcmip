netcdf CFS-atmos-northPacific-Pair-1995 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:36:53 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1995/roms-cfs-atmos-Pair-1995.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1995/CFS-atmos-northPacific-Pair-1995.nc\n",
			"Mon Sep 10 13:31:31 2018: Time overhang added\n",
			"Mon Sep 10 13:31:27 2018: ncrcat /tmp/tpcdf23897_6d7e_43be_9af4_ad293bf03618.nc frc/roms-cfs-atmos-Pair-1995.nc /tmp/tpb84e6d01_15f2_4aa0_9e51_b0b9bfd4ce96.nc /tmp/tpdde4c4ed_fb03_451c_9eca_7334f183619b.nc\n",
			"Mon Sep 10 13:31:27 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-1995.nc /tmp/tpcdf23897_6d7e_43be_9af4_ad293bf03618.nc\n",
			"Thu Sep  6 09:49:33 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1995.nc\n",
			"Thu Sep  6 09:48:35 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_1995_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-1995.nc\n",
			"04-Oct-2017 17:36:52: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
