netcdf CFS-atmos-northPacific-Vwind-2013 {
dimensions:
	wind_time = UNLIMITED ; // (1448 currently)
	lat = 342 ;
	lon = 587 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:23:07 2022: ncks -F -O -d wind_time,2,1449 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2013/roms-cfs-atmos-Vwind-2013.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2013/CFS-atmos-northPacific-Vwind-2013.nc\n",
			"Mon Sep 10 13:45:27 2018: Time overhang added\n",
			"Mon Sep 10 13:45:19 2018: ncrcat /tmp/tpd86b60a3_139f_49da_aa81_0b5bfa7d8db1.nc frc/roms-cfs-atmos-Vwind-2013.nc /tmp/tp96dac500_4252_4b1d_8c9a_7f862af1698d.nc /tmp/tp928f0fe4_19bd_4cf8_b386_2fde4d4c0de1.nc\n",
			"Mon Sep 10 13:45:19 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2013.nc /tmp/tpd86b60a3_139f_49da_aa81_0b5bfa7d8db1.nc\n",
			"Thu Sep  6 13:09:07 2018: ncks -O -F -d wind_time,2,1449 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2013_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2013.nc\n",
			"04-Oct-2017 18:23:31: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
