netcdf CFS-ocean-ESPER-Bering10K-N30-brycarbon-2007 {
dimensions:
	bry_time = UNLIMITED ; // (73 currently)
	s_rho = 30 ;
	eta_rho = 258 ;
	xi_rho = 182 ;
variables:
	double bry_time(bry_time) ;
		bry_time:long_name = "time since initialization" ;
		bry_time:units = "seconds since 1900-01-01 00:00:00" ;
		bry_time:calendar = "standard" ;
		bry_time:cell_methods = "bry_time: mean" ;
	double salt_east(bry_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity, eastern boundary condition" ;
		salt_east:time = "bry_time" ;
		salt_east:cell_methods = "bry_time: mean" ;
	double salt_south(bry_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity, southern boundary condition" ;
		salt_south:time = "bry_time" ;
		salt_south:cell_methods = "bry_time: mean" ;
	double salt_west(bry_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity, western boundary condition" ;
		salt_west:time = "bry_time" ;
		salt_west:cell_methods = "bry_time: mean" ;
	double alkalinity_west(bry_time, s_rho, eta_rho) ;
		alkalinity_west:long_name = "alkalinity western boundary condition" ;
		alkalinity_west:units = "umol/kg" ;
		alkalinity_west:time = "bry_time" ;
		alkalinity_west:_FillValue = 1.e+36 ;
	double TIC_west(bry_time, s_rho, eta_rho) ;
		TIC_west:long_name = "TIC western boundary condition" ;
		TIC_west:units = "umol/kg" ;
		TIC_west:time = "bry_time" ;
		TIC_west:_FillValue = 1.e+36 ;
	double alkalinity_east(bry_time, s_rho, eta_rho) ;
		alkalinity_east:long_name = "alkalinity eastern boundary condition" ;
		alkalinity_east:units = "umol/kg" ;
		alkalinity_east:time = "bry_time" ;
		alkalinity_east:_FillValue = 1.e+36 ;
	double TIC_east(bry_time, s_rho, eta_rho) ;
		TIC_east:long_name = "TIC eastern boundary condition" ;
		TIC_east:units = "umol/kg" ;
		TIC_east:time = "bry_time" ;
		TIC_east:_FillValue = 1.e+36 ;
	double alkalinity_south(bry_time, s_rho, xi_rho) ;
		alkalinity_south:long_name = "alkalinity southern boundary condition" ;
		alkalinity_south:units = "umol/kg" ;
		alkalinity_south:time = "bry_time" ;
		alkalinity_south:_FillValue = 1.e+36 ;
	double TIC_south(bry_time, s_rho, xi_rho) ;
		TIC_south:long_name = "TIC southern boundary condition" ;
		TIC_south:units = "umol/kg" ;
		TIC_south:time = "bry_time" ;
		TIC_south:_FillValue = 1.e+36 ;

// global attributes:
		:type = "BOUNDARY file" ;
		:history = "Tue Jan 17 15:49:37 2023: TIC and alkalinity estimated by salinty regression via ESPER_Mixed\n",
			"Tue Jan 17 15:48:00 2023: ncks -v salt_west,salt_east,salt_south /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2007/CFS-ocean-Bering10K-N30-bryocn-2007.nc /Users/kakearney/Documents/Research/Working/mox_bumblereem/ROMS_Datasets/CFS/2007/CFS-ocean-ESPER-Bering10K-N30-brycarbon-2007.nc\n",
			"Tue Dec 27 21:26:32 2022: ncrcat -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad02.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad03.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad04.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad05.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad06.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad07.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad08.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad09.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad10.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad11.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad12.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad13.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad14.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad15.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad16.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad17.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad18.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad19.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad20.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad21.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad22.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad23.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad24.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad25.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad26.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad27.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad28.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad29.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad30.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad31.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad32.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad33.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad34.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad35.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad36.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad37.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad38.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad39.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad40.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad41.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad42.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad43.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad44.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad45.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad46.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad47.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad48.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad49.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad50.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad51.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad52.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad53.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad54.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad55.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad56.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad57.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad58.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad59.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad60.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad61.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad62.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad63.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad64.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad65.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad66.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad67.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad68.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad69.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad70.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad71.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad72.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad73.nc <>/final/2007/CFS-ocean-Bering10K-N30-bryocn-2007.nc\n",
			"Tue Dec 27 21:25:10 2022: ncks -O -F -d s_rho,1,30 <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad01.nc\n",
			"Tue Dec 27 21:25:09 2022: ncra -O <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad01.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad01.nc\n",
			"Tue Dec 27 21:25:09 2022: ncrcat -O <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010100.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010106.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010112.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010118.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010200.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010206.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010212.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010218.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010300.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010306.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010312.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010318.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010400.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010406.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010412.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010418.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010500.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010506.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010512.nc <>/prep/singletime/CFS-ocean-Bering10K-N30-bryocn-2007010518.nc <>/prep/pentads/CFS-ocean-Bering10K-N30-bryocn-2007pentad01.nc\n",
			"Tue Dec 27 06:39:23 2022: CFS data added\n",
			"Tue Dec 20 15:09:11 2022: File schema created via bry_schema.m" ;
		:NCO = "netCDF Operators version 5.1.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
