netcdf CFS-atmos-northPacific-Pair-2018 {
dimensions:
	pair_time = UNLIMITED ; // (1452 currently)
	lat = 344 ;
	lon = 588 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:missing_value = -1.e+34 ;
		Pair:_FillValue = -1.e+34 ;
		Pair:time = "pair_time" ;
		Pair:coordinates = "lon lat" ;
		Pair:long_name = "atmos pressure" ;
		Pair:history = "From roms-cfs-atmos-Pair-2018" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double pair_time(pair_time) ;
		pair_time:units = "day since 1900-01-01 00:00:00" ;
		pair_time:time_origin = "01-JAN-1900 00:00:00" ;
		pair_time:axis = "T" ;
		pair_time:standard_name = "time" ;

// global attributes:
		:history = "Mon Oct 31 12:21:41 2022: ncks -F -O -d pair_time,2,1453 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Pair-2018.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2018/CFS-atmos-northPacific-Pair-2018.nc\n",
			"Thu May 30 20:48:31 2019: Time overhang added\n",
			"Thu May 30 20:48:24 2019: ncrcat /tmp/tpbe60aebc_cc7b_4dde_92a3_25d2afedbd87.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Pair-2018.nc /tmp/tp50601ae6_4161_4240_a236_d2888e42b47d.nc /tmp/tp4d3dfef6_f975_4505_9514_aacba959955a.nc\n",
			"Thu May 30 20:48:23 2019: ncks -F -d pair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2018/roms-cfs-atmos-Pair-2018.nc /tmp/tpbe60aebc_cc7b_4dde_92a3_25d2afedbd87.nc\n",
			"FERRET V7.4  29-May-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
