netcdf CFS-atmos-northPacific-Pair-1984 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 225 ;
	lon = 385 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:missing_value = -1.e+34 ;
		Pair:_FillValue = -1.e+34 ;
		Pair:time = "pair_time" ;
		Pair:coordinates = "lon lat" ;
		Pair:long_name = "atmos pressure" ;
		Pair:history = "From roms-cfs-atmos-Pair-1984" ;
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double pair_time(pair_time) ;
		pair_time:units = "day since 1900-01-01 00:00:00" ;
		pair_time:time_origin = "01-JAN-1900 00:00:00" ;
		pair_time:axis = "T" ;
		pair_time:standard_name = "time" ;

// global attributes:
		:history = "Thu Nov  3 15:34:18 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Pair-1984.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1984/CFS-atmos-northPacific-Pair-1984.nc\n",
			"Wed Nov 20 13:43:58 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:43:54 2019: ncrcat /tmp/tpad15a540_7a03_47d1_945a_6bd22f2efaf1.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Pair-1984.nc /tmp/tpfe6534bc_4788_48cc_9f63_d8dd40a70cf3.nc /tmp/tpd9862338_abf0_4e35_bdce_a9869f33f114.nc\n",
			"Wed Nov 20 13:43:52 2019: ncks -F -d pair_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-Pair-1984.nc /tmp/tpad15a540_7a03_47d1_945a_6bd22f2efaf1.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
