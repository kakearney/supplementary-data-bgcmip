netcdf CFS-atmos-northPacific-Vwind-2005 {
dimensions:
	wind_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Vwind(wind_time, lat, lon) ;
		Vwind:long_name = "surface v-wind component" ;
		Vwind:units = "meter second-1" ;
		Vwind:coordinates = "lon lat" ;
		Vwind:time = "wind_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double wind_time(wind_time) ;
		wind_time:long_name = "forcing time" ;
		wind_time:units = "days since 1900-01-01 00:00:00" ;
		wind_time:time = "wind_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:51:52 2022: ncks -F -O -d wind_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2005/roms-cfs-atmos-Vwind-2005.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2005/CFS-atmos-northPacific-Vwind-2005.nc\n",
			"Mon Sep 10 13:44:24 2018: Time overhang added\n",
			"Mon Sep 10 13:44:20 2018: ncrcat /tmp/tpc4165d69_ff37_46fd_baf4_80e7801fe32b.nc frc/roms-cfs-atmos-Vwind-2005.nc /tmp/tped2c6f5a_6d44_43a2_a79f_67068c72a4f5.nc /tmp/tp3fd54905_5d5d_41ff_a53d_0057a63ca13b.nc\n",
			"Mon Sep 10 13:44:20 2018: ncks -F -d wind_time,1,1 frc/roms-cfs-atmos-Vwind-2005.nc /tmp/tpc4165d69_ff37_46fd_baf4_80e7801fe32b.nc\n",
			"Thu Sep  6 11:24:44 2018: ncks -O -F -d wind_time,2,1461 -v Vwind /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2005_wind.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Vwind-2005.nc\n",
			"04-Oct-2017 18:02:37: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
