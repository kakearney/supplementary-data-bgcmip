netcdf CFS-atmos-northPacific-rain-2011 {
dimensions:
	lat = 342 ;
	lon = 587 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double rain(rain_time, lat, lon) ;
		rain:long_name = "rain fall rate" ;
		rain:units = "kilogram meter-2 second-1" ;
		rain:coordinates = "lon lat" ;
		rain:time = "rain_time" ;
	double rain_time(rain_time) ;
		rain_time:long_name = "forcing time" ;
		rain_time:units = "days since 1900-01-01 00:00:00" ;
		rain_time:time = "rain_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 17:12:32 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2011/roms-cfs-atmos-rain-2011.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2011/CFS-atmos-northPacific-rain-2011.nc\n",
			"Mon Sep 10 13:51:26 2018: Time overhang added\n",
			"Mon Sep 10 13:51:18 2018: ncrcat /tmp/tp733d5d56_2fca_4293_9d12_79e9c5d5033f.nc frc/roms-cfs-atmos-rain-2011.nc /tmp/tpfa40d3ed_82f9_4c9e_afcd_bf2e52b20c94.nc /tmp/tp4959d8a2_7ecd_45e9_aab9_4fbb1cbf6fd6.nc\n",
			"Mon Sep 10 13:51:17 2018: ncks -F -d rain_time,1,1 frc/roms-cfs-atmos-rain-2011.nc /tmp/tp733d5d56_2fca_4293_9d12_79e9c5d5033f.nc\n",
			"Thu Sep  6 12:27:15 2018: ncks -O -F -d rain_time,2,1461 /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2011_rain.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-rain-2011.nc\n",
			"04-Oct-2017 18:16:43: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
