netcdf CFS-atmos-northPacific-rain-1984 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	rain_time = UNLIMITED ; // (1460 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double rain(rain_time, lat, lon) ;
		rain:missing_value = -1.e+34 ;
		rain:_FillValue = -1.e+34 ;
		rain:time = "rain_time" ;
		rain:coordinates = "lon lat" ;
		rain:long_name = "rainfall" ;
		rain:history = "From roms-cfs-atmos-rain-1984" ;
	double rain_time(rain_time) ;
		rain_time:units = "day since 1900-01-01 00:00:00" ;
		rain_time:time_origin = "01-JAN-1900 00:00:00" ;
		rain_time:axis = "T" ;
		rain_time:standard_name = "time" ;

// global attributes:
		:history = "Thu Nov  3 15:35:12 2022: ncks -F -O -d rain_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-rain-1984.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1984/CFS-atmos-northPacific-rain-1984.nc\n",
			"Wed Nov 20 13:45:25 2019: Time overhang added to both ends\n",
			"Wed Nov 20 13:45:18 2019: ncrcat /tmp/tpb7c119f3_bf90_41c2_8a18_19f13d7bc6eb.nc /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-rain-1984.nc /tmp/tp814f4f6c_73fc_42df_9e0e_73e7126b6ffc.nc /tmp/tp9e5330ca_cf7d_43ad_92f1_c87a57484fb0.nc\n",
			"Wed Nov 20 13:45:16 2019: ncks -F -d rain_time,1,1 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1984/roms-cfs-atmos-rain-1984.nc /tmp/tpb7c119f3_bf90_41c2_8a18_19f13d7bc6eb.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
