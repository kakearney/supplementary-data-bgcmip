netcdf CFS-atmos-northPacific-rain-1985 {
dimensions:
	lat = 225 ;
	lon = 385 ;
	rain_time = UNLIMITED ; // (1459 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:point_spacing = "uneven" ;
		lat:axis = "Y" ;
		lat:standard_name = "latitude" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:modulo = 360.f ;
		lon:point_spacing = "uneven" ;
		lon:axis = "X" ;
		lon:standard_name = "longitude" ;
	double rain(rain_time, lat, lon) ;
		rain:missing_value = -1.e+34 ;
		rain:_FillValue = -1.e+34 ;
		rain:time = "rain_time" ;
		rain:coordinates = "lon lat" ;
		rain:long_name = "rainfall" ;
		rain:history = "From roms-cfs-atmos-rain-1985" ;
	double rain_time(rain_time) ;
		rain_time:units = "day since 1900-01-01 00:00:00" ;
		rain_time:time_origin = "01-JAN-1900 00:00:00" ;
		rain_time:axis = "T" ;
		rain_time:standard_name = "time" ;

// global attributes:
		:history = "Fri Oct 28 16:19:16 2022: ncks -F -O -d rain_time,2,1460 /gscratch/bumblereem/bering10k/input/hindcast_cfs/1985/roms-cfs-atmos-rain-1985.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/1985/CFS-atmos-northPacific-rain-1985.nc\n",
			"Wed Nov 20 13:47:22 2019: Time overhang added to end\n",
			"Wed Nov 20 13:47:18 2019: ncrcat /gscratch/bumblereem/bering10k/input/hindcast_cfs/1985/roms-cfs-atmos-rain-1985.nc /tmp/tp75b9b11d_b907_4701_8bb2_1407d3bb72ea.nc /tmp/tp48414017_eda1_4d9f_ab76_1ba71c9f3d18.nc\n",
			"FERRET V7.4  11-Oct-19" ;
		:Conventions = "CF-1.6" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
