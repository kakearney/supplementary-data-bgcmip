netcdf CFS-atmos-northPacific-Pair-2003 {
dimensions:
	pair_time = UNLIMITED ; // (1460 currently)
	lat = 224 ;
	lon = 384 ;
variables:
	double Pair(pair_time, lat, lon) ;
		Pair:long_name = "surface air pressure" ;
		Pair:units = "Pascal" ;
		Pair:coordinates = "lon lat" ;
		Pair:time = "air_time" ;
	double lat(lat, lon) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:coordinates = "lon lat" ;
	double lon(lat, lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:coordinates = "lon lat" ;
	double pair_time(pair_time) ;
		pair_time:long_name = "forcing time" ;
		pair_time:units = "days since 1900-01-01 00:00:00" ;
		pair_time:time = "air_time" ;

// global attributes:
		:type = "FORCING file" ;
		:title = "Hindcast surface flux forcing for Bering 10K ROMS domain" ;
		:history = "Fri Oct 28 16:16:50 2022: ncks -F -O -d pair_time,2,1461 /gscratch/bumblereem/bering10k/input/hindcast_cfs/2003/roms-cfs-atmos-Pair-2003.nc /gscratch/bumblereem/kearney/ROMS_Datasets/CFS/2003/CFS-atmos-northPacific-Pair-2003.nc\n",
			"Mon Sep 10 13:32:23 2018: Time overhang added\n",
			"Mon Sep 10 13:32:19 2018: ncrcat /tmp/tpc9c37e9d_7712_40f2_bc3a_a8b46ac2b838.nc frc/roms-cfs-atmos-Pair-2003.nc /tmp/tp81d6a563_18ce_4097_b039_043c3a648a52.nc /tmp/tpa33069ff_bf4d_405d_8908_28a588265a0a.nc\n",
			"Mon Sep 10 13:32:19 2018: ncks -F -d pair_time,1,1 frc/roms-cfs-atmos-Pair-2003.nc /tmp/tpc9c37e9d_7712_40f2_bc3a_a8b46ac2b838.nc\n",
			"Thu Sep  6 10:59:59 2018: ncrename -d air_time,pair_time -v air_time,pair_time /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2003.nc\n",
			"Thu Sep  6 10:58:53 2018: ncks -O -F -d air_time,2,1461 -v Pair /Volumes/Storage/BeringROMS/hindcastFrcBry/frc/corecfs_2003_air.nc /Volumes/Storage/BeringROMS/hindcastFrcBry/CFS/roms-cfs-atmos-Pair-2003.nc\n",
			"04-Oct-2017 17:57:09: File schema defined via bering10k_schema.m" ;
		:NCO = "4.6.9" ;
		:nco_openmp_thread_number = 1 ;
}
